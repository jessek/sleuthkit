<!doctype html><html lang="en-US" dir="ltr"><head><base href="https://accounts.google.com/v3/signin/"><link rel="preconnect" href="//www.gstatic.com"><meta name="referrer" content="origin"><style data-href="https://www.gstatic.com/_/mss/boq-identity/_/ss/k=boq-identity.AccountsSignInUi.V77lomOXnCU.L.W.O/am=iQEMSyZrAIVyBAAUAgBAAIACAAAAAAAAAEBgAACACQE/d=1/ed=1/rs=AOaEmlEhiUj1HQAWI5Xn5Zignm3WIbgnLA/m=identifierview,_b,_tp" nonce="D3in5SeEvI-f7-RWiq5EjQ">@-webkit-keyframes quantumWizBoxInkSpread{0%{-webkit-transform:translate(-50%,-50%) scale(0.2);-webkit-transform:translate(-50%,-50%) scale(0.2);transform:translate(-50%,-50%) scale(0.2)}to{-webkit-transform:translate(-50%,-50%) scale(2.2);-webkit-transform:translate(-50%,-50%) scale(2.2);transform:translate(-50%,-50%) scale(2.2)}}@keyframes quantumWizBoxInkSpread{0%{-webkit-transform:translate(-50%,-50%) scale(0.2);-webkit-transform:translate(-50%,-50%) scale(0.2);transform:translate(-50%,-50%) scale(0.2)}to{-webkit-transform:translate(-50%,-50%) scale(2.2);-webkit-transform:translate(-50%,-50%) scale(2.2);transform:translate(-50%,-50%) scale(2.2)}}@-webkit-keyframes quantumWizIconFocusPulse{0%{-webkit-transform:translate(-50%,-50%) scale(1.5);-webkit-transform:translate(-50%,-50%) scale(1.5);transform:translate(-50%,-50%) scale(1.5);opacity:0}to{-webkit-transform:translate(-50%,-50%) scale(2);-webkit-transform:translate(-50%,-50%) scale(2);transform:translate(-50%,-50%) scale(2);opacity:1}}@keyframes quantumWizIconFocusPulse{0%{-webkit-transform:translate(-50%,-50%) scale(1.5);-webkit-transform:translate(-50%,-50%) scale(1.5);transform:translate(-50%,-50%) scale(1.5);opacity:0}to{-webkit-transform:translate(-50%,-50%) scale(2);-webkit-transform:translate(-50%,-50%) scale(2);transform:translate(-50%,-50%) scale(2);opacity:1}}@-webkit-keyframes quantumWizRadialInkSpread{0%{-webkit-transform:scale(1.5);-webkit-transform:scale(1.5);transform:scale(1.5);opacity:0}to{-webkit-transform:scale(2.5);-webkit-transform:scale(2.5);transform:scale(2.5);opacity:1}}@keyframes quantumWizRadialInkSpread{0%{-webkit-transform:scale(1.5);-webkit-transform:scale(1.5);transform:scale(1.5);opacity:0}to{-webkit-transform:scale(2.5);-webkit-transform:scale(2.5);transform:scale(2.5);opacity:1}}@-webkit-keyframes quantumWizRadialInkFocusPulse{0%{-webkit-transform:scale(2);-webkit-transform:scale(2);transform:scale(2);opacity:0}to{-webkit-transform:scale(2.5);-webkit-transform:scale(2.5);transform:scale(2.5);opacity:1}}@keyframes quantumWizRadialInkFocusPulse{0%{-webkit-transform:scale(2);-webkit-transform:scale(2);transform:scale(2);opacity:0}to{-webkit-transform:scale(2.5);-webkit-transform:scale(2.5);transform:scale(2.5);opacity:1}}@-webkit-keyframes mdc-ripple-fg-radius-in{0%{-webkit-animation-timing-function:cubic-bezier(0.4,0,0.2,1);-webkit-animation-timing-function:cubic-bezier(0.4,0,0.2,1);animation-timing-function:cubic-bezier(0.4,0,0.2,1);-webkit-transform:translate(var(--mdc-ripple-fg-translate-start,0)) scale(1);-webkit-transform:translate(var(--mdc-ripple-fg-translate-start,0)) scale(1);transform:translate(var(--mdc-ripple-fg-translate-start,0)) scale(1)}to{-webkit-transform:translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1));-webkit-transform:translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1));transform:translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1))}}@keyframes mdc-ripple-fg-radius-in{0%{-webkit-animation-timing-function:cubic-bezier(0.4,0,0.2,1);-webkit-animation-timing-function:cubic-bezier(0.4,0,0.2,1);animation-timing-function:cubic-bezier(0.4,0,0.2,1);-webkit-transform:translate(var(--mdc-ripple-fg-translate-start,0)) scale(1);-webkit-transform:translate(var(--mdc-ripple-fg-translate-start,0)) scale(1);transform:translate(var(--mdc-ripple-fg-translate-start,0)) scale(1)}to{-webkit-transform:translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1));-webkit-transform:translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1));transform:translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1))}}@-webkit-keyframes mdc-ripple-fg-opacity-in{0%{-webkit-animation-timing-function:linear;-webkit-animation-timing-function:linear;animation-timing-function:linear;opacity:0}to{opacity:var(--mdc-ripple-fg-opacity,0)}}@keyframes mdc-ripple-fg-opacity-in{0%{-webkit-animation-timing-function:linear;-webkit-animation-timing-function:linear;animation-timing-function:linear;opacity:0}to{opacity:var(--mdc-ripple-fg-opacity,0)}}@-webkit-keyframes mdc-ripple-fg-opacity-out{0%{-webkit-animation-timing-function:linear;-webkit-animation-timing-function:linear;animation-timing-function:linear;opacity:var(--mdc-ripple-fg-opacity,0)}to{opacity:0}}@keyframes mdc-ripple-fg-opacity-out{0%{-webkit-animation-timing-function:linear;-webkit-animation-timing-function:linear;animation-timing-function:linear;opacity:var(--mdc-ripple-fg-opacity,0)}to{opacity:0}}.VfPpkd-ksKsZd-XxIAqe{--mdc-ripple-fg-size:0;--mdc-ripple-left:0;--mdc-ripple-top:0;--mdc-ripple-fg-scale:1;--mdc-ripple-fg-translate-end:0;--mdc-ripple-fg-translate-start:0;-webkit-tap-highlight-color:rgba(0,0,0,0);will-change:transform,opacity;position:relative;outline:none;overflow:hidden}.VfPpkd-ksKsZd-XxIAqe::before,.VfPpkd-ksKsZd-XxIAqe::after{position:absolute;-webkit-border-radius:50%;border-radius:50%;opacity:0;pointer-events:none;content:""}.VfPpkd-ksKsZd-XxIAqe::before{-webkit-transition:opacity 15ms linear,background-color 15ms linear;-webkit-transition:opacity 15ms linear,background-color 15ms linear;transition:opacity 15ms linear,background-color 15ms linear;z-index:1;z-index:var(--mdc-ripple-z-index,1)}.VfPpkd-ksKsZd-XxIAqe::after{z-index:0;z-index:var(--mdc-ripple-z-index,0)}.VfPpkd-ksKsZd-XxIAqe.VfPpkd-ksKsZd-mWPk3d::before{-webkit-transform:scale(var(--mdc-ripple-fg-scale,1));-webkit-transform:scale(var(--mdc-ripple-fg-scale,1));transform:scale(var(--mdc-ripple-fg-scale,1))}.VfPpkd-ksKsZd-XxIAqe.VfPpkd-ksKsZd-mWPk3d::after{top:0;left:0;-webkit-transform:scale(0);-webkit-transform:scale(0);transform:scale(0);-webkit-transform-origin:center center;-webkit-transform-origin:center center;transform-origin:center center}.VfPpkd-ksKsZd-XxIAqe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd::after{top:var(--mdc-ripple-top,0);left:var(--mdc-ripple-left,0)}.VfPpkd-ksKsZd-XxIAqe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-lJfZMc::after{-webkit-animation:mdc-ripple-fg-radius-in 225ms forwards,mdc-ripple-fg-opacity-in 75ms forwards;-webkit-animation:mdc-ripple-fg-radius-in 225ms forwards,mdc-ripple-fg-opacity-in 75ms forwards;animation:mdc-ripple-fg-radius-in 225ms forwards,mdc-ripple-fg-opacity-in 75ms forwards}.VfPpkd-ksKsZd-XxIAqe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-OmS1vf::after{-webkit-animation:mdc-ripple-fg-opacity-out 150ms;-webkit-animation:mdc-ripple-fg-opacity-out 150ms;animation:mdc-ripple-fg-opacity-out 150ms;-webkit-transform:translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1));-webkit-transform:translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1));transform:translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1))}.VfPpkd-ksKsZd-XxIAqe::before,.VfPpkd-ksKsZd-XxIAqe::after{top:-webkit-calc(50% - 100%);top:calc(50% - 100%);left:-webkit-calc(50% - 100%);left:calc(50% - 100%);width:200%;height:200%}.VfPpkd-ksKsZd-XxIAqe.VfPpkd-ksKsZd-mWPk3d::after{width:var(--mdc-ripple-fg-size,100%);height:var(--mdc-ripple-fg-size,100%)}.VfPpkd-ksKsZd-XxIAqe[data-mdc-ripple-is-unbounded],.VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd{overflow:visible}.VfPpkd-ksKsZd-XxIAqe[data-mdc-ripple-is-unbounded]::before,.VfPpkd-ksKsZd-XxIAqe[data-mdc-ripple-is-unbounded]::after,.VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd::before,.VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd::after{top:-webkit-calc(50% - 50%);top:calc(50% - 50%);left:-webkit-calc(50% - 50%);left:calc(50% - 50%);width:100%;height:100%}.VfPpkd-ksKsZd-XxIAqe[data-mdc-ripple-is-unbounded].VfPpkd-ksKsZd-mWPk3d::before,.VfPpkd-ksKsZd-XxIAqe[data-mdc-ripple-is-unbounded].VfPpkd-ksKsZd-mWPk3d::after,.VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd.VfPpkd-ksKsZd-mWPk3d::before,.VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd.VfPpkd-ksKsZd-mWPk3d::after{top:var(--mdc-ripple-top,calc(50% - 50%));left:var(--mdc-ripple-left,calc(50% - 50%));width:var(--mdc-ripple-fg-size,100%);height:var(--mdc-ripple-fg-size,100%)}.VfPpkd-ksKsZd-XxIAqe[data-mdc-ripple-is-unbounded].VfPpkd-ksKsZd-mWPk3d::after,.VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd.VfPpkd-ksKsZd-mWPk3d::after{width:var(--mdc-ripple-fg-size,100%);height:var(--mdc-ripple-fg-size,100%)}.VfPpkd-ksKsZd-XxIAqe::before,.VfPpkd-ksKsZd-XxIAqe::after{background-color:#000;background-color:var(--mdc-ripple-color,#000)}.VfPpkd-ksKsZd-XxIAqe:hover::before,.VfPpkd-ksKsZd-XxIAqe.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,0.04)}.VfPpkd-ksKsZd-XxIAqe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe::before,.VfPpkd-ksKsZd-XxIAqe:not(.VfPpkd-ksKsZd-mWPk3d):focus::before{-webkit-transition-duration:75ms;-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,0.12)}.VfPpkd-ksKsZd-XxIAqe:not(.VfPpkd-ksKsZd-mWPk3d)::after{-webkit-transition:opacity 150ms linear;-webkit-transition:opacity 150ms linear;transition:opacity 150ms linear}.VfPpkd-ksKsZd-XxIAqe:not(.VfPpkd-ksKsZd-mWPk3d):active::after{-webkit-transition-duration:75ms;-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-press-opacity,0.12)}.VfPpkd-ksKsZd-XxIAqe.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.12)}.VfPpkd-Bz112c-LgbsSe{font-size:24px;width:48px;height:48px;padding:12px}.VfPpkd-Bz112c-LgbsSe.VfPpkd-Bz112c-LgbsSe-OWXEXe-e5LLRc-SxQuSe .VfPpkd-Bz112c-Jh9lGc{width:40px;height:40px;margin-top:4px;margin-bottom:4px;margin-right:4px;margin-left:4px}.VfPpkd-Bz112c-LgbsSe.VfPpkd-Bz112c-LgbsSe-OWXEXe-e5LLRc-SxQuSe .VfPpkd-Bz112c-J1Ukfc-LhBDec{max-height:40px;max-width:40px}.VfPpkd-Bz112c-LgbsSe:disabled{color:rgba(0,0,0,.38);color:var(--mdc-theme-text-disabled-on-light,rgba(0,0,0,.38))}.VfPpkd-Bz112c-LgbsSe svg,.VfPpkd-Bz112c-LgbsSe img{width:24px;height:24px}.VfPpkd-Bz112c-LgbsSe{display:inline-block;position:relative;box-sizing:border-box;border:none;outline:none;background-color:transparent;fill:currentColor;color:inherit;text-decoration:none;cursor:pointer;-webkit-user-select:none;user-select:none;z-index:0;overflow:visible}.VfPpkd-Bz112c-LgbsSe .VfPpkd-Bz112c-RLmnJb{position:absolute;top:50%;height:48px;left:50%;width:48px;-webkit-transform:translate(-50%,-50%);transform:translate(-50%,-50%)}@media screen and (forced-colors:active){.VfPpkd-Bz112c-LgbsSe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Bz112c-J1Ukfc-LhBDec,.VfPpkd-Bz112c-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Bz112c-J1Ukfc-LhBDec{display:block}}.VfPpkd-Bz112c-LgbsSe:disabled{cursor:default;pointer-events:none}.VfPpkd-Bz112c-LgbsSe[hidden]{display:none}.VfPpkd-Bz112c-LgbsSe-OWXEXe-KVuj8d-Q3DXx{-webkit-box-align:center;-webkit-align-items:center;align-items:center;display:-webkit-inline-box;display:-webkit-inline-flex;display:inline-flex;-webkit-box-pack:center;-webkit-justify-content:center;justify-content:center}.VfPpkd-Bz112c-J1Ukfc-LhBDec{pointer-events:none;border:2px solid transparent;border-radius:6px;box-sizing:content-box;position:absolute;top:50%;left:50%;-webkit-transform:translate(-50%,-50%);transform:translate(-50%,-50%);height:100%;width:100%;display:none}@media screen and (forced-colors:active){.VfPpkd-Bz112c-J1Ukfc-LhBDec{border-color:CanvasText}}.VfPpkd-Bz112c-J1Ukfc-LhBDec::after{content:"";border:2px solid transparent;border-radius:8px;display:block;position:absolute;top:50%;left:50%;-webkit-transform:translate(-50%,-50%);transform:translate(-50%,-50%);height:calc(100% + 4px);width:calc(100% + 4px)}@media screen and (forced-colors:active){.VfPpkd-Bz112c-J1Ukfc-LhBDec::after{border-color:CanvasText}}.VfPpkd-Bz112c-kBDsod{display:inline-block}.VfPpkd-Bz112c-kBDsod.VfPpkd-Bz112c-kBDsod-OWXEXe-IT5dJd,.VfPpkd-Bz112c-LgbsSe-OWXEXe-IT5dJd .VfPpkd-Bz112c-kBDsod{display:none}.VfPpkd-Bz112c-LgbsSe-OWXEXe-IT5dJd .VfPpkd-Bz112c-kBDsod.VfPpkd-Bz112c-kBDsod-OWXEXe-IT5dJd{display:inline-block}.VfPpkd-Bz112c-mRLv6{height:100%;left:0;outline:none;position:absolute;top:0;width:100%}.VfPpkd-Bz112c-LgbsSe{--mdc-ripple-fg-size:0;--mdc-ripple-left:0;--mdc-ripple-top:0;--mdc-ripple-fg-scale:1;--mdc-ripple-fg-translate-end:0;--mdc-ripple-fg-translate-start:0;-webkit-tap-highlight-color:rgba(0,0,0,0);will-change:transform,opacity}.VfPpkd-Bz112c-LgbsSe .VfPpkd-Bz112c-Jh9lGc::before,.VfPpkd-Bz112c-LgbsSe .VfPpkd-Bz112c-Jh9lGc::after{position:absolute;border-radius:50%;opacity:0;pointer-events:none;content:""}.VfPpkd-Bz112c-LgbsSe .VfPpkd-Bz112c-Jh9lGc::before{-webkit-transition:opacity 15ms linear,background-color 15ms linear;transition:opacity 15ms linear,background-color 15ms linear;z-index:1;z-index:var(--mdc-ripple-z-index,1)}.VfPpkd-Bz112c-LgbsSe .VfPpkd-Bz112c-Jh9lGc::after{z-index:0;z-index:var(--mdc-ripple-z-index,0)}.VfPpkd-Bz112c-LgbsSe.VfPpkd-ksKsZd-mWPk3d .VfPpkd-Bz112c-Jh9lGc::before{-webkit-transform:scale(var(--mdc-ripple-fg-scale,1));transform:scale(var(--mdc-ripple-fg-scale,1))}.VfPpkd-Bz112c-LgbsSe.VfPpkd-ksKsZd-mWPk3d .VfPpkd-Bz112c-Jh9lGc::after{top:0;left:0;-webkit-transform:scale(0);transform:scale(0);-webkit-transform-origin:center center;transform-origin:center center}.VfPpkd-Bz112c-LgbsSe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd .VfPpkd-Bz112c-Jh9lGc::after{top:var(--mdc-ripple-top,0);left:var(--mdc-ripple-left,0)}.VfPpkd-Bz112c-LgbsSe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-lJfZMc .VfPpkd-Bz112c-Jh9lGc::after{-webkit-animation:mdc-ripple-fg-radius-in 225ms forwards,mdc-ripple-fg-opacity-in 75ms forwards;animation:mdc-ripple-fg-radius-in 225ms forwards,mdc-ripple-fg-opacity-in 75ms forwards}.VfPpkd-Bz112c-LgbsSe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-OmS1vf .VfPpkd-Bz112c-Jh9lGc::after{-webkit-animation:mdc-ripple-fg-opacity-out .15s;animation:mdc-ripple-fg-opacity-out .15s;-webkit-transform:translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1));transform:translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1))}.VfPpkd-Bz112c-LgbsSe .VfPpkd-Bz112c-Jh9lGc::before,.VfPpkd-Bz112c-LgbsSe .VfPpkd-Bz112c-Jh9lGc::after{top:0;left:0;width:100%;height:100%}.VfPpkd-Bz112c-LgbsSe.VfPpkd-ksKsZd-mWPk3d .VfPpkd-Bz112c-Jh9lGc::before,.VfPpkd-Bz112c-LgbsSe.VfPpkd-ksKsZd-mWPk3d .VfPpkd-Bz112c-Jh9lGc::after{top:var(--mdc-ripple-top,0);left:var(--mdc-ripple-left,0);width:var(--mdc-ripple-fg-size,100%);height:var(--mdc-ripple-fg-size,100%)}.VfPpkd-Bz112c-LgbsSe.VfPpkd-ksKsZd-mWPk3d .VfPpkd-Bz112c-Jh9lGc::after{width:var(--mdc-ripple-fg-size,100%);height:var(--mdc-ripple-fg-size,100%)}.VfPpkd-Bz112c-LgbsSe .VfPpkd-Bz112c-Jh9lGc::before,.VfPpkd-Bz112c-LgbsSe .VfPpkd-Bz112c-Jh9lGc::after{background-color:#000;background-color:var(--mdc-ripple-color,#000)}.VfPpkd-Bz112c-LgbsSe:hover .VfPpkd-Bz112c-Jh9lGc::before,.VfPpkd-Bz112c-LgbsSe.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Bz112c-Jh9lGc::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.VfPpkd-Bz112c-LgbsSe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Bz112c-Jh9lGc::before,.VfPpkd-Bz112c-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Bz112c-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.VfPpkd-Bz112c-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Bz112c-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.VfPpkd-Bz112c-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Bz112c-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-press-opacity,.12)}.VfPpkd-Bz112c-LgbsSe.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.12)}.VfPpkd-Bz112c-LgbsSe:disabled:hover .VfPpkd-Bz112c-Jh9lGc::before,.VfPpkd-Bz112c-LgbsSe:disabled.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Bz112c-Jh9lGc::before{opacity:0;opacity:var(--mdc-ripple-hover-opacity,0)}.VfPpkd-Bz112c-LgbsSe:disabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Bz112c-Jh9lGc::before,.VfPpkd-Bz112c-LgbsSe:disabled:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Bz112c-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:0;opacity:var(--mdc-ripple-focus-opacity,0)}.VfPpkd-Bz112c-LgbsSe:disabled:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Bz112c-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.VfPpkd-Bz112c-LgbsSe:disabled:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Bz112c-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:0;opacity:var(--mdc-ripple-press-opacity,0)}.VfPpkd-Bz112c-LgbsSe:disabled.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0)}.VfPpkd-Bz112c-LgbsSe .VfPpkd-Bz112c-Jh9lGc{height:100%;left:0;pointer-events:none;position:absolute;top:0;width:100%;z-index:-1}.VfPpkd-dgl2Hf-ppHlrf-sM5MNb{display:inline}.VfPpkd-LgbsSe{position:relative;display:-webkit-inline-box;display:-webkit-inline-flex;display:inline-flex;-webkit-box-align:center;-webkit-align-items:center;align-items:center;-webkit-box-pack:center;-webkit-justify-content:center;justify-content:center;box-sizing:border-box;min-width:64px;border:none;outline:none;line-height:inherit;-webkit-user-select:none;user-select:none;-webkit-appearance:none;overflow:visible;vertical-align:middle;background:transparent}.VfPpkd-LgbsSe .VfPpkd-BFbNVe-bF1uUb{width:100%;height:100%;top:0;left:0}.VfPpkd-LgbsSe::-moz-focus-inner{padding:0;border:0}.VfPpkd-LgbsSe:active{outline:none}.VfPpkd-LgbsSe:hover{cursor:pointer}.VfPpkd-LgbsSe:disabled{cursor:default;pointer-events:none}.VfPpkd-LgbsSe[hidden]{display:none}.VfPpkd-LgbsSe .VfPpkd-kBDsod{margin-left:0;margin-right:8px;display:inline-block;position:relative;vertical-align:top}[dir=rtl] .VfPpkd-LgbsSe .VfPpkd-kBDsod,.VfPpkd-LgbsSe .VfPpkd-kBDsod[dir=rtl]{margin-left:8px;margin-right:0}.VfPpkd-LgbsSe .VfPpkd-UdE5de-uDEFge{font-size:0;position:absolute;-webkit-transform:translate(-50%,-50%);transform:translate(-50%,-50%);top:50%;left:50%;line-height:normal}.VfPpkd-LgbsSe .VfPpkd-vQzf8d{position:relative}.VfPpkd-LgbsSe .VfPpkd-J1Ukfc-LhBDec{pointer-events:none;border:2px solid transparent;border-radius:6px;box-sizing:content-box;position:absolute;top:50%;left:50%;-webkit-transform:translate(-50%,-50%);transform:translate(-50%,-50%);height:calc(100% + 4px);width:calc(100% + 4px);display:none}@media screen and (forced-colors:active){.VfPpkd-LgbsSe .VfPpkd-J1Ukfc-LhBDec{border-color:CanvasText}}.VfPpkd-LgbsSe .VfPpkd-J1Ukfc-LhBDec::after{content:"";border:2px solid transparent;border-radius:8px;display:block;position:absolute;top:50%;left:50%;-webkit-transform:translate(-50%,-50%);transform:translate(-50%,-50%);height:calc(100% + 4px);width:calc(100% + 4px)}@media screen and (forced-colors:active){.VfPpkd-LgbsSe .VfPpkd-J1Ukfc-LhBDec::after{border-color:CanvasText}}@media screen and (forced-colors:active){.VfPpkd-LgbsSe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-J1Ukfc-LhBDec,.VfPpkd-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-J1Ukfc-LhBDec{display:block}}.VfPpkd-LgbsSe .VfPpkd-RLmnJb{position:absolute;top:50%;height:48px;left:0;right:0;-webkit-transform:translateY(-50%);transform:translateY(-50%)}.VfPpkd-vQzf8d+.VfPpkd-kBDsod{margin-left:8px;margin-right:0}[dir=rtl] .VfPpkd-vQzf8d+.VfPpkd-kBDsod,.VfPpkd-vQzf8d+.VfPpkd-kBDsod[dir=rtl]{margin-left:0;margin-right:8px}svg.VfPpkd-kBDsod{fill:currentColor}.VfPpkd-LgbsSe-OWXEXe-dgl2Hf{margin-top:6px;margin-bottom:6px}.VfPpkd-LgbsSe{-moz-osx-font-smoothing:grayscale;-webkit-font-smoothing:antialiased;text-decoration:none}.VfPpkd-LgbsSe{padding:0 8px 0 8px}.VfPpkd-LgbsSe-OWXEXe-k8QpJ{-webkit-transition:box-shadow .28s cubic-bezier(.4,0,.2,1);transition:box-shadow .28s cubic-bezier(.4,0,.2,1);padding:0 16px 0 16px}.VfPpkd-LgbsSe-OWXEXe-k8QpJ.VfPpkd-LgbsSe-OWXEXe-Bz112c-UbuQg{padding:0 12px 0 16px}.VfPpkd-LgbsSe-OWXEXe-k8QpJ.VfPpkd-LgbsSe-OWXEXe-Bz112c-M1Soyc{padding:0 16px 0 12px}.VfPpkd-LgbsSe-OWXEXe-MV7yeb{-webkit-transition:box-shadow .28s cubic-bezier(.4,0,.2,1);transition:box-shadow .28s cubic-bezier(.4,0,.2,1);padding:0 16px 0 16px}.VfPpkd-LgbsSe-OWXEXe-MV7yeb.VfPpkd-LgbsSe-OWXEXe-Bz112c-UbuQg{padding:0 12px 0 16px}.VfPpkd-LgbsSe-OWXEXe-MV7yeb.VfPpkd-LgbsSe-OWXEXe-Bz112c-M1Soyc{padding:0 16px 0 12px}.VfPpkd-LgbsSe-OWXEXe-INsAgc{border-style:solid;-webkit-transition:border .28s cubic-bezier(.4,0,.2,1);transition:border .28s cubic-bezier(.4,0,.2,1)}.VfPpkd-LgbsSe-OWXEXe-INsAgc .VfPpkd-Jh9lGc{border-style:solid;border-color:transparent}.VfPpkd-LgbsSe{--mdc-ripple-fg-size:0;--mdc-ripple-left:0;--mdc-ripple-top:0;--mdc-ripple-fg-scale:1;--mdc-ripple-fg-translate-end:0;--mdc-ripple-fg-translate-start:0;-webkit-tap-highlight-color:rgba(0,0,0,0);will-change:transform,opacity}.VfPpkd-LgbsSe .VfPpkd-Jh9lGc::before,.VfPpkd-LgbsSe .VfPpkd-Jh9lGc::after{position:absolute;border-radius:50%;opacity:0;pointer-events:none;content:""}.VfPpkd-LgbsSe .VfPpkd-Jh9lGc::before{-webkit-transition:opacity 15ms linear,background-color 15ms linear;transition:opacity 15ms linear,background-color 15ms linear;z-index:1}.VfPpkd-LgbsSe .VfPpkd-Jh9lGc::after{z-index:0}.VfPpkd-LgbsSe.VfPpkd-ksKsZd-mWPk3d .VfPpkd-Jh9lGc::before{-webkit-transform:scale(var(--mdc-ripple-fg-scale,1));transform:scale(var(--mdc-ripple-fg-scale,1))}.VfPpkd-LgbsSe.VfPpkd-ksKsZd-mWPk3d .VfPpkd-Jh9lGc::after{top:0;left:0;-webkit-transform:scale(0);transform:scale(0);-webkit-transform-origin:center center;transform-origin:center center}.VfPpkd-LgbsSe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd .VfPpkd-Jh9lGc::after{top:var(--mdc-ripple-top,0);left:var(--mdc-ripple-left,0)}.VfPpkd-LgbsSe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-lJfZMc .VfPpkd-Jh9lGc::after{-webkit-animation:mdc-ripple-fg-radius-in 225ms forwards,mdc-ripple-fg-opacity-in 75ms forwards;animation:mdc-ripple-fg-radius-in 225ms forwards,mdc-ripple-fg-opacity-in 75ms forwards}.VfPpkd-LgbsSe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-OmS1vf .VfPpkd-Jh9lGc::after{-webkit-animation:mdc-ripple-fg-opacity-out .15s;animation:mdc-ripple-fg-opacity-out .15s;-webkit-transform:translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1));transform:translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1))}.VfPpkd-LgbsSe .VfPpkd-Jh9lGc::before,.VfPpkd-LgbsSe .VfPpkd-Jh9lGc::after{top:-50%;left:-50%;width:200%;height:200%}.VfPpkd-LgbsSe.VfPpkd-ksKsZd-mWPk3d .VfPpkd-Jh9lGc::after{width:var(--mdc-ripple-fg-size,100%);height:var(--mdc-ripple-fg-size,100%)}.VfPpkd-Jh9lGc{position:absolute;box-sizing:content-box;overflow:hidden;z-index:0;top:0;left:0;bottom:0;right:0}.VfPpkd-LgbsSe{font-family:Roboto,sans-serif;font-size:.875rem;letter-spacing:.0892857143em;font-weight:500;text-transform:uppercase;height:36px;border-radius:4px}.VfPpkd-LgbsSe:not(:disabled){color:#6200ee}.VfPpkd-LgbsSe:disabled{color:rgba(0,0,0,.38)}.VfPpkd-LgbsSe .VfPpkd-kBDsod{font-size:1.125rem;width:1.125rem;height:1.125rem}.VfPpkd-LgbsSe .VfPpkd-Jh9lGc::before{background-color:#6200ee}.VfPpkd-LgbsSe .VfPpkd-Jh9lGc::after{background-color:#6200ee}.VfPpkd-LgbsSe:hover .VfPpkd-Jh9lGc::before,.VfPpkd-LgbsSe.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:.04}.VfPpkd-LgbsSe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.VfPpkd-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12}.VfPpkd-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.VfPpkd-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12}.VfPpkd-LgbsSe.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-text-button-pressed-state-layer-opacity,0.12)}.VfPpkd-LgbsSe .VfPpkd-Jh9lGc{border-radius:4px}.VfPpkd-LgbsSe .VfPpkd-J1Ukfc-LhBDec{border-radius:2px}.VfPpkd-LgbsSe .VfPpkd-J1Ukfc-LhBDec::after{border-radius:4px}.VfPpkd-LgbsSe-OWXEXe-k8QpJ{font-family:Roboto,sans-serif;font-size:.875rem;letter-spacing:.0892857143em;font-weight:500;text-transform:uppercase;height:36px;border-radius:4px}.VfPpkd-LgbsSe-OWXEXe-k8QpJ:not(:disabled){background-color:#6200ee}.VfPpkd-LgbsSe-OWXEXe-k8QpJ:disabled{background-color:rgba(0,0,0,.12)}.VfPpkd-LgbsSe-OWXEXe-k8QpJ:not(:disabled){color:#fff}.VfPpkd-LgbsSe-OWXEXe-k8QpJ:disabled{color:rgba(0,0,0,.38)}.VfPpkd-LgbsSe-OWXEXe-k8QpJ .VfPpkd-kBDsod{font-size:1.125rem;width:1.125rem;height:1.125rem}.VfPpkd-LgbsSe-OWXEXe-k8QpJ .VfPpkd-Jh9lGc::before{background-color:#fff}.VfPpkd-LgbsSe-OWXEXe-k8QpJ .VfPpkd-Jh9lGc::after{background-color:#fff}.VfPpkd-LgbsSe-OWXEXe-k8QpJ:hover .VfPpkd-Jh9lGc::before,.VfPpkd-LgbsSe-OWXEXe-k8QpJ.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:.08}.VfPpkd-LgbsSe-OWXEXe-k8QpJ.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.VfPpkd-LgbsSe-OWXEXe-k8QpJ:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.24}.VfPpkd-LgbsSe-OWXEXe-k8QpJ:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.VfPpkd-LgbsSe-OWXEXe-k8QpJ:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.24}.VfPpkd-LgbsSe-OWXEXe-k8QpJ.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-filled-button-pressed-state-layer-opacity,0.24)}.VfPpkd-LgbsSe-OWXEXe-k8QpJ .VfPpkd-Jh9lGc{border-radius:4px}.VfPpkd-LgbsSe-OWXEXe-k8QpJ .VfPpkd-J1Ukfc-LhBDec{border-radius:2px}.VfPpkd-LgbsSe-OWXEXe-k8QpJ .VfPpkd-J1Ukfc-LhBDec::after{border-radius:4px}.VfPpkd-LgbsSe-OWXEXe-MV7yeb{font-family:Roboto,sans-serif;font-size:.875rem;letter-spacing:.0892857143em;font-weight:500;text-transform:uppercase;height:36px;border-radius:4px;box-shadow:0 3px 1px -2px rgba(0,0,0,.2),0 2px 2px 0 rgba(0,0,0,.14),0 1px 5px 0 rgba(0,0,0,.12)}.VfPpkd-LgbsSe-OWXEXe-MV7yeb:not(:disabled){background-color:#6200ee}.VfPpkd-LgbsSe-OWXEXe-MV7yeb:disabled{background-color:rgba(0,0,0,.12)}.VfPpkd-LgbsSe-OWXEXe-MV7yeb:not(:disabled){color:#fff}.VfPpkd-LgbsSe-OWXEXe-MV7yeb:disabled{color:rgba(0,0,0,.38)}.VfPpkd-LgbsSe-OWXEXe-MV7yeb .VfPpkd-kBDsod{font-size:1.125rem;width:1.125rem;height:1.125rem}.VfPpkd-LgbsSe-OWXEXe-MV7yeb .VfPpkd-Jh9lGc::before{background-color:#fff}.VfPpkd-LgbsSe-OWXEXe-MV7yeb .VfPpkd-Jh9lGc::after{background-color:#fff}.VfPpkd-LgbsSe-OWXEXe-MV7yeb:hover .VfPpkd-Jh9lGc::before,.VfPpkd-LgbsSe-OWXEXe-MV7yeb.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:.08}.VfPpkd-LgbsSe-OWXEXe-MV7yeb.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.VfPpkd-LgbsSe-OWXEXe-MV7yeb:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.24}.VfPpkd-LgbsSe-OWXEXe-MV7yeb:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.VfPpkd-LgbsSe-OWXEXe-MV7yeb:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.24}.VfPpkd-LgbsSe-OWXEXe-MV7yeb.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-protected-button-pressed-state-layer-opacity,0.24)}.VfPpkd-LgbsSe-OWXEXe-MV7yeb .VfPpkd-Jh9lGc{border-radius:4px}.VfPpkd-LgbsSe-OWXEXe-MV7yeb .VfPpkd-J1Ukfc-LhBDec{border-radius:2px}.VfPpkd-LgbsSe-OWXEXe-MV7yeb .VfPpkd-J1Ukfc-LhBDec::after{border-radius:4px}.VfPpkd-LgbsSe-OWXEXe-MV7yeb.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.VfPpkd-LgbsSe-OWXEXe-MV7yeb:not(.VfPpkd-ksKsZd-mWPk3d):focus{box-shadow:0 2px 4px -1px rgba(0,0,0,.2),0 4px 5px 0 rgba(0,0,0,.14),0 1px 10px 0 rgba(0,0,0,.12)}.VfPpkd-LgbsSe-OWXEXe-MV7yeb:hover{box-shadow:0 2px 4px -1px rgba(0,0,0,.2),0 4px 5px 0 rgba(0,0,0,.14),0 1px 10px 0 rgba(0,0,0,.12)}.VfPpkd-LgbsSe-OWXEXe-MV7yeb:not(:disabled):active{box-shadow:0 5px 5px -3px rgba(0,0,0,.2),0 8px 10px 1px rgba(0,0,0,.14),0 3px 14px 2px rgba(0,0,0,.12)}.VfPpkd-LgbsSe-OWXEXe-MV7yeb:disabled{box-shadow:0 0 0 0 rgba(0,0,0,.2),0 0 0 0 rgba(0,0,0,.14),0 0 0 0 rgba(0,0,0,.12)}.VfPpkd-LgbsSe-OWXEXe-INsAgc{font-family:Roboto,sans-serif;font-size:.875rem;letter-spacing:.0892857143em;font-weight:500;text-transform:uppercase;height:36px;border-radius:4px;padding:0 15px 0 15px;border-width:1px}.VfPpkd-LgbsSe-OWXEXe-INsAgc:not(:disabled){color:#6200ee}.VfPpkd-LgbsSe-OWXEXe-INsAgc:disabled{color:rgba(0,0,0,.38)}.VfPpkd-LgbsSe-OWXEXe-INsAgc .VfPpkd-kBDsod{font-size:1.125rem;width:1.125rem;height:1.125rem}.VfPpkd-LgbsSe-OWXEXe-INsAgc .VfPpkd-Jh9lGc::before{background-color:#6200ee}.VfPpkd-LgbsSe-OWXEXe-INsAgc .VfPpkd-Jh9lGc::after{background-color:#6200ee}.VfPpkd-LgbsSe-OWXEXe-INsAgc:hover .VfPpkd-Jh9lGc::before,.VfPpkd-LgbsSe-OWXEXe-INsAgc.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:.04}.VfPpkd-LgbsSe-OWXEXe-INsAgc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.VfPpkd-LgbsSe-OWXEXe-INsAgc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12}.VfPpkd-LgbsSe-OWXEXe-INsAgc:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.VfPpkd-LgbsSe-OWXEXe-INsAgc:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12}.VfPpkd-LgbsSe-OWXEXe-INsAgc.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-outlined-button-pressed-state-layer-opacity,0.12)}.VfPpkd-LgbsSe-OWXEXe-INsAgc .VfPpkd-Jh9lGc{border-radius:4px}.VfPpkd-LgbsSe-OWXEXe-INsAgc .VfPpkd-J1Ukfc-LhBDec{border-radius:2px}.VfPpkd-LgbsSe-OWXEXe-INsAgc .VfPpkd-J1Ukfc-LhBDec::after{border-radius:4px}.VfPpkd-LgbsSe-OWXEXe-INsAgc:not(:disabled){border-color:rgba(0,0,0,.12)}.VfPpkd-LgbsSe-OWXEXe-INsAgc:disabled{border-color:rgba(0,0,0,.12)}.VfPpkd-LgbsSe-OWXEXe-INsAgc.VfPpkd-LgbsSe-OWXEXe-Bz112c-UbuQg{padding:0 11px 0 15px}.VfPpkd-LgbsSe-OWXEXe-INsAgc.VfPpkd-LgbsSe-OWXEXe-Bz112c-M1Soyc{padding:0 15px 0 11px}.VfPpkd-LgbsSe-OWXEXe-INsAgc .VfPpkd-Jh9lGc{top:-1px;left:-1px;bottom:-1px;right:-1px;border-width:1px}.VfPpkd-LgbsSe-OWXEXe-INsAgc .VfPpkd-RLmnJb{left:-1px;width:calc(100% + 2px)}.nCP5yc{font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:.875rem;letter-spacing:.0107142857em;font-weight:500;text-transform:none;-webkit-transition:border .28s cubic-bezier(.4,0,.2,1),box-shadow .28s cubic-bezier(.4,0,.2,1);transition:border .28s cubic-bezier(.4,0,.2,1),box-shadow .28s cubic-bezier(.4,0,.2,1);box-shadow:none}.nCP5yc .VfPpkd-Jh9lGc{height:100%;position:absolute;overflow:hidden;width:100%;z-index:0}.nCP5yc:not(:disabled){background-color:rgb(26,115,232);background-color:var(--gm-fillbutton-container-color,rgb(26,115,232))}.nCP5yc:not(:disabled){color:#fff;color:var(--gm-fillbutton-ink-color,#fff)}.nCP5yc:disabled{background-color:rgba(60,64,67,.12);background-color:var(--gm-fillbutton-disabled-container-color,rgba(60,64,67,.12))}.nCP5yc:disabled{color:rgba(60,64,67,.38);color:var(--gm-fillbutton-disabled-ink-color,rgba(60,64,67,.38))}.nCP5yc .VfPpkd-Jh9lGc::before,.nCP5yc .VfPpkd-Jh9lGc::after{background-color:rgb(32,33,36);background-color:var(--gm-fillbutton-state-color,rgb(32,33,36))}.nCP5yc:hover .VfPpkd-Jh9lGc::before,.nCP5yc.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:.16;opacity:var(--mdc-ripple-hover-opacity,.16)}.nCP5yc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.nCP5yc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.24;opacity:var(--mdc-ripple-focus-opacity,.24)}.nCP5yc:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.nCP5yc:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.2;opacity:var(--mdc-ripple-press-opacity,.2)}.nCP5yc.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.2)}.nCP5yc .VfPpkd-BFbNVe-bF1uUb{opacity:0}.nCP5yc .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo,.nCP5yc .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:#fff}@media (-ms-high-contrast:active),screen and (forced-colors:active){.nCP5yc .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo,.nCP5yc .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:CanvasText}}.nCP5yc:hover{box-shadow:0 1px 2px 0 rgba(60,64,67,.3),0 1px 3px 1px rgba(60,64,67,.15);box-shadow:0 1px 2px 0 var(--gm-fillbutton-keyshadow-color,rgba(60,64,67,.3)),0 1px 3px 1px var(--gm-fillbutton-ambientshadow-color,rgba(60,64,67,.15))}.nCP5yc:hover .VfPpkd-BFbNVe-bF1uUb{opacity:0}.nCP5yc:active{box-shadow:0 1px 2px 0 rgba(60,64,67,.3),0 2px 6px 2px rgba(60,64,67,.15);box-shadow:0 1px 2px 0 var(--gm-fillbutton-keyshadow-color,rgba(60,64,67,.3)),0 2px 6px 2px var(--gm-fillbutton-ambientshadow-color,rgba(60,64,67,.15))}.nCP5yc:active .VfPpkd-BFbNVe-bF1uUb{opacity:0}.nCP5yc:disabled{box-shadow:none}.nCP5yc:disabled:hover .VfPpkd-Jh9lGc::before,.nCP5yc:disabled.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:0;opacity:var(--mdc-ripple-hover-opacity,0)}.nCP5yc:disabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.nCP5yc:disabled:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:0;opacity:var(--mdc-ripple-focus-opacity,0)}.nCP5yc:disabled:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.nCP5yc:disabled:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:0;opacity:var(--mdc-ripple-press-opacity,0)}.nCP5yc:disabled.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0)}.nCP5yc:disabled .VfPpkd-BFbNVe-bF1uUb{opacity:0}.Rj2Mlf{font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:.875rem;letter-spacing:.0107142857em;font-weight:500;text-transform:none;-webkit-transition:border .28s cubic-bezier(.4,0,.2,1),box-shadow .28s cubic-bezier(.4,0,.2,1);transition:border .28s cubic-bezier(.4,0,.2,1),box-shadow .28s cubic-bezier(.4,0,.2,1);box-shadow:none}.Rj2Mlf .VfPpkd-Jh9lGc{height:100%;position:absolute;overflow:hidden;width:100%;z-index:0}.Rj2Mlf:not(:disabled){color:rgb(26,115,232);color:var(--gm-hairlinebutton-ink-color,rgb(26,115,232))}.Rj2Mlf:not(:disabled){border-color:rgb(218,220,224);border-color:var(--gm-hairlinebutton-outline-color,rgb(218,220,224))}.Rj2Mlf:not(:disabled):hover{border-color:rgb(218,220,224);border-color:var(--gm-hairlinebutton-outline-color,rgb(218,220,224))}.Rj2Mlf:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.Rj2Mlf:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{border-color:rgb(23,78,166);border-color:var(--gm-hairlinebutton-outline-color--stateful,rgb(23,78,166))}.Rj2Mlf:not(:disabled):active,.Rj2Mlf:not(:disabled):focus:active{border-color:rgb(218,220,224);border-color:var(--gm-hairlinebutton-outline-color,rgb(218,220,224))}.Rj2Mlf:disabled{color:rgba(60,64,67,.38);color:var(--gm-hairlinebutton-disabled-ink-color,rgba(60,64,67,.38))}.Rj2Mlf:disabled{border-color:rgba(60,64,67,.12);border-color:var(--gm-hairlinebutton-disabled-outline-color,rgba(60,64,67,.12))}.Rj2Mlf:hover:not(:disabled),.Rj2Mlf.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:disabled),.Rj2Mlf:not(.VfPpkd-ksKsZd-mWPk3d):focus:not(:disabled),.Rj2Mlf:active:not(:disabled){color:rgb(23,78,166);color:var(--gm-hairlinebutton-ink-color--stateful,rgb(23,78,166))}.Rj2Mlf .VfPpkd-BFbNVe-bF1uUb{opacity:0}.Rj2Mlf .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo,.Rj2Mlf .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:rgb(26,115,232)}@media (-ms-high-contrast:active),screen and (forced-colors:active){.Rj2Mlf .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo,.Rj2Mlf .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:CanvasText}}.Rj2Mlf .VfPpkd-Jh9lGc::before,.Rj2Mlf .VfPpkd-Jh9lGc::after{background-color:rgb(26,115,232);background-color:var(--gm-hairlinebutton-state-color,rgb(26,115,232))}.Rj2Mlf:hover .VfPpkd-Jh9lGc::before,.Rj2Mlf.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.Rj2Mlf.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.Rj2Mlf:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.Rj2Mlf:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.Rj2Mlf:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-press-opacity,.12)}.Rj2Mlf.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.12)}.Rj2Mlf:disabled:hover .VfPpkd-Jh9lGc::before,.Rj2Mlf:disabled.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:0;opacity:var(--mdc-ripple-hover-opacity,0)}.Rj2Mlf:disabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.Rj2Mlf:disabled:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:0;opacity:var(--mdc-ripple-focus-opacity,0)}.Rj2Mlf:disabled:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.Rj2Mlf:disabled:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:0;opacity:var(--mdc-ripple-press-opacity,0)}.Rj2Mlf:disabled.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0)}.b9hyVd{font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:.875rem;letter-spacing:.0107142857em;font-weight:500;text-transform:none;-webkit-transition:border .28s cubic-bezier(.4,0,.2,1),box-shadow .28s cubic-bezier(.4,0,.2,1);transition:border .28s cubic-bezier(.4,0,.2,1),box-shadow .28s cubic-bezier(.4,0,.2,1);border-width:0;box-shadow:0 1px 2px 0 rgba(60,64,67,.3),0 1px 3px 1px rgba(60,64,67,.15);box-shadow:0 1px 2px 0 var(--gm-protectedbutton-keyshadow-color,rgba(60,64,67,.3)),0 1px 3px 1px var(--gm-protectedbutton-ambientshadow-color,rgba(60,64,67,.15))}.b9hyVd .VfPpkd-Jh9lGc{height:100%;position:absolute;overflow:hidden;width:100%;z-index:0}.b9hyVd:not(:disabled){background-color:#fff;background-color:var(--gm-protectedbutton-container-color,#fff)}.b9hyVd:not(:disabled){color:rgb(26,115,232);color:var(--gm-protectedbutton-ink-color,rgb(26,115,232))}.b9hyVd:disabled{background-color:rgba(60,64,67,.12);background-color:var(--gm-protectedbutton-disabled-container-color,rgba(60,64,67,.12))}.b9hyVd:disabled{color:rgba(60,64,67,.38);color:var(--gm-protectedbutton-disabled-ink-color,rgba(60,64,67,.38))}.b9hyVd:hover:not(:disabled),.b9hyVd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:disabled),.b9hyVd:not(.VfPpkd-ksKsZd-mWPk3d):focus:not(:disabled),.b9hyVd:active:not(:disabled){color:rgb(23,78,166);color:var(--gm-protectedbutton-ink-color--stateful,rgb(23,78,166))}.b9hyVd .VfPpkd-BFbNVe-bF1uUb{opacity:0}.b9hyVd .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo,.b9hyVd .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:rgb(26,115,232)}@media (-ms-high-contrast:active),screen and (forced-colors:active){.b9hyVd .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo,.b9hyVd .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:CanvasText}}.b9hyVd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.b9hyVd:not(.VfPpkd-ksKsZd-mWPk3d):focus{border-width:0;box-shadow:0 1px 2px 0 rgba(60,64,67,.3),0 1px 3px 1px rgba(60,64,67,.15);box-shadow:0 1px 2px 0 var(--gm-protectedbutton-keyshadow-color,rgba(60,64,67,.3)),0 1px 3px 1px var(--gm-protectedbutton-ambientshadow-color,rgba(60,64,67,.15))}.b9hyVd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-BFbNVe-bF1uUb,.b9hyVd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-BFbNVe-bF1uUb{opacity:0}.b9hyVd:hover{border-width:0;box-shadow:0 1px 2px 0 rgba(60,64,67,.3),0 2px 6px 2px rgba(60,64,67,.15);box-shadow:0 1px 2px 0 var(--gm-protectedbutton-keyshadow-color,rgba(60,64,67,.3)),0 2px 6px 2px var(--gm-protectedbutton-ambientshadow-color,rgba(60,64,67,.15))}.b9hyVd:hover .VfPpkd-BFbNVe-bF1uUb{opacity:0}.b9hyVd:not(:disabled):active{border-width:0;box-shadow:0 1px 3px 0 rgba(60,64,67,.3),0 4px 8px 3px rgba(60,64,67,.15);box-shadow:0 1px 3px 0 var(--gm-protectedbutton-keyshadow-color,rgba(60,64,67,.3)),0 4px 8px 3px var(--gm-protectedbutton-ambientshadow-color,rgba(60,64,67,.15))}.b9hyVd:not(:disabled):active .VfPpkd-BFbNVe-bF1uUb{opacity:0}.b9hyVd .VfPpkd-Jh9lGc::before,.b9hyVd .VfPpkd-Jh9lGc::after{background-color:rgb(26,115,232);background-color:var(--gm-protectedbutton-state-color,rgb(26,115,232))}.b9hyVd:hover .VfPpkd-Jh9lGc::before,.b9hyVd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.b9hyVd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.b9hyVd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.b9hyVd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.b9hyVd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-press-opacity,.12)}.b9hyVd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.12)}.b9hyVd:disabled{box-shadow:none}.b9hyVd:disabled .VfPpkd-BFbNVe-bF1uUb{opacity:0}.b9hyVd:disabled:hover .VfPpkd-Jh9lGc::before,.b9hyVd:disabled.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:0;opacity:var(--mdc-ripple-hover-opacity,0)}.b9hyVd:disabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.b9hyVd:disabled:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:0;opacity:var(--mdc-ripple-focus-opacity,0)}.b9hyVd:disabled:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.b9hyVd:disabled:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:0;opacity:var(--mdc-ripple-press-opacity,0)}.b9hyVd:disabled.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0)}.Kjnxrf{font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:.875rem;letter-spacing:.0107142857em;font-weight:500;text-transform:none;-webkit-transition:border .28s cubic-bezier(.4,0,.2,1),box-shadow .28s cubic-bezier(.4,0,.2,1);transition:border .28s cubic-bezier(.4,0,.2,1),box-shadow .28s cubic-bezier(.4,0,.2,1);box-shadow:none}.Kjnxrf .VfPpkd-Jh9lGc{height:100%;position:absolute;overflow:hidden;width:100%;z-index:0}.Kjnxrf:not(:disabled){background-color:rgb(232,240,254)}.Kjnxrf:not(:disabled){color:rgb(25,103,210)}.Kjnxrf:disabled{background-color:rgba(60,64,67,.12)}.Kjnxrf:disabled{color:rgba(60,64,67,.38)}.Kjnxrf:hover:not(:disabled),.Kjnxrf.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:disabled),.Kjnxrf:not(.VfPpkd-ksKsZd-mWPk3d):focus:not(:disabled),.Kjnxrf:active:not(:disabled){color:rgb(23,78,166)}.Kjnxrf .VfPpkd-Jh9lGc::before,.Kjnxrf .VfPpkd-Jh9lGc::after{background-color:rgb(25,103,210);background-color:var(--mdc-ripple-color,rgb(25,103,210))}.Kjnxrf:hover .VfPpkd-Jh9lGc::before,.Kjnxrf.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.Kjnxrf.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.Kjnxrf:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.Kjnxrf:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.Kjnxrf:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.Kjnxrf.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}.Kjnxrf .VfPpkd-BFbNVe-bF1uUb{opacity:0}.Kjnxrf .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo,.Kjnxrf .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:rgb(25,103,210)}@media (-ms-high-contrast:active),screen and (forced-colors:active){.Kjnxrf .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo,.Kjnxrf .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:CanvasText}}.Kjnxrf:hover{box-shadow:0 1px 2px 0 rgba(60,64,67,.3),0 1px 3px 1px rgba(60,64,67,.15)}.Kjnxrf:hover .VfPpkd-BFbNVe-bF1uUb{opacity:0}.Kjnxrf:not(:disabled):active{box-shadow:0 1px 2px 0 rgba(60,64,67,.3),0 2px 6px 2px rgba(60,64,67,.15)}.Kjnxrf:not(:disabled):active .VfPpkd-BFbNVe-bF1uUb{opacity:0}.Kjnxrf:disabled{box-shadow:none}.Kjnxrf:disabled .VfPpkd-BFbNVe-bF1uUb{opacity:0}.Kjnxrf:disabled:hover .VfPpkd-Jh9lGc::before,.Kjnxrf:disabled.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:0;opacity:var(--mdc-ripple-hover-opacity,0)}.Kjnxrf:disabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.Kjnxrf:disabled:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:0;opacity:var(--mdc-ripple-focus-opacity,0)}.Kjnxrf:disabled:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.Kjnxrf:disabled:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:0;opacity:var(--mdc-ripple-press-opacity,0)}.Kjnxrf:disabled.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0)}.ksBjEc{font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:.875rem;letter-spacing:.0107142857em;font-weight:500;text-transform:none}.ksBjEc .VfPpkd-Jh9lGc{height:100%;position:absolute;overflow:hidden;width:100%;z-index:0}.ksBjEc:not(:disabled){background-color:transparent}.ksBjEc:not(:disabled){color:rgb(26,115,232);color:var(--gm-colortextbutton-ink-color,rgb(26,115,232))}.ksBjEc:disabled{color:rgba(60,64,67,.38);color:var(--gm-colortextbutton-disabled-ink-color,rgba(60,64,67,.38))}.ksBjEc .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo,.ksBjEc .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:rgb(26,115,232)}@media (-ms-high-contrast:active),screen and (forced-colors:active){.ksBjEc .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo,.ksBjEc .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:CanvasText}}.ksBjEc:hover:not(:disabled),.ksBjEc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:disabled),.ksBjEc:not(.VfPpkd-ksKsZd-mWPk3d):focus:not(:disabled),.ksBjEc:active:not(:disabled){color:rgb(23,78,166);color:var(--gm-colortextbutton-ink-color--stateful,rgb(23,78,166))}.ksBjEc .VfPpkd-Jh9lGc::before,.ksBjEc .VfPpkd-Jh9lGc::after{background-color:rgb(26,115,232);background-color:var(--gm-colortextbutton-state-color,rgb(26,115,232))}.ksBjEc:hover .VfPpkd-Jh9lGc::before,.ksBjEc.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.ksBjEc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.ksBjEc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.ksBjEc:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.ksBjEc:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-press-opacity,.12)}.ksBjEc.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.12)}.ksBjEc:disabled:hover .VfPpkd-Jh9lGc::before,.ksBjEc:disabled.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:0;opacity:var(--mdc-ripple-hover-opacity,0)}.ksBjEc:disabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.ksBjEc:disabled:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:0;opacity:var(--mdc-ripple-focus-opacity,0)}.ksBjEc:disabled:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.ksBjEc:disabled:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:0;opacity:var(--mdc-ripple-press-opacity,0)}.ksBjEc:disabled.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0)}.LjDxcd{font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:.875rem;letter-spacing:.0107142857em;font-weight:500;text-transform:none}.LjDxcd .VfPpkd-Jh9lGc{height:100%;position:absolute;overflow:hidden;width:100%;z-index:0}.LjDxcd:not(:disabled){color:rgb(95,99,104);color:var(--gm-neutraltextbutton-ink-color,rgb(95,99,104))}.LjDxcd:disabled{color:rgba(60,64,67,.38);color:var(--gm-neutraltextbutton-disabled-ink-color,rgba(60,64,67,.38))}.LjDxcd:hover:not(:disabled),.LjDxcd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:disabled),.LjDxcd:not(.VfPpkd-ksKsZd-mWPk3d):focus:not(:disabled),.LjDxcd:active:not(:disabled){color:rgb(32,33,36);color:var(--gm-neutraltextbutton-ink-color--stateful,rgb(32,33,36))}.LjDxcd .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo,.LjDxcd .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:rgb(95,99,104)}@media (-ms-high-contrast:active),screen and (forced-colors:active){.LjDxcd .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo,.LjDxcd .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:CanvasText}}.LjDxcd .VfPpkd-Jh9lGc::before,.LjDxcd .VfPpkd-Jh9lGc::after{background-color:rgb(95,99,104);background-color:var(--gm-neutraltextbutton-state-color,rgb(95,99,104))}.LjDxcd:hover .VfPpkd-Jh9lGc::before,.LjDxcd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.LjDxcd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.LjDxcd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.LjDxcd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.LjDxcd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-press-opacity,.12)}.LjDxcd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.12)}.LjDxcd:disabled:hover .VfPpkd-Jh9lGc::before,.LjDxcd:disabled.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:0;opacity:var(--mdc-ripple-hover-opacity,0)}.LjDxcd:disabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.LjDxcd:disabled:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:0;opacity:var(--mdc-ripple-focus-opacity,0)}.LjDxcd:disabled:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.LjDxcd:disabled:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:0;opacity:var(--mdc-ripple-press-opacity,0)}.LjDxcd:disabled.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0)}.DuMIQc{padding:0 24px 0 24px}.P62QJc{padding:0 23px 0 23px;border-width:1px}.P62QJc.VfPpkd-LgbsSe-OWXEXe-Bz112c-UbuQg{padding:0 11px 0 23px}.P62QJc.VfPpkd-LgbsSe-OWXEXe-Bz112c-M1Soyc{padding:0 23px 0 11px}.P62QJc .VfPpkd-Jh9lGc{top:-1px;left:-1px;bottom:-1px;right:-1px;border-width:1px}.P62QJc .VfPpkd-RLmnJb{left:-1px;width:calc(100% + 2px)}.yHy1rc{z-index:0}.yHy1rc .VfPpkd-Bz112c-Jh9lGc::before,.yHy1rc .VfPpkd-Bz112c-Jh9lGc::after{z-index:-1}.yHy1rc:disabled{color:rgba(60,64,67,.38);color:var(--gm-iconbutton-disabled-ink-color,rgba(60,64,67,.38))}.fzRBVc{z-index:0}.fzRBVc .VfPpkd-Bz112c-Jh9lGc::before,.fzRBVc .VfPpkd-Bz112c-Jh9lGc::after{z-index:-1}.fzRBVc:disabled{color:rgba(60,64,67,.38);color:var(--gm-iconbutton-disabled-ink-color,rgba(60,64,67,.38))}.WpHeLc{height:100%;left:0;position:absolute;top:0;width:100%;outline:none}[dir=rtl] .HDnnrf .VfPpkd-kBDsod,.HDnnrf .VfPpkd-kBDsod[dir=rtl]{-webkit-transform:scaleX(-1);transform:scaleX(-1)}[dir=rtl] .QDwDD,.QDwDD[dir=rtl]{-webkit-transform:scaleX(-1);transform:scaleX(-1)}.PDpWxe{will-change:unset}.LQeN7 .VfPpkd-J1Ukfc-LhBDec{pointer-events:none;border:2px solid rgb(24,90,188);border-radius:6px;box-sizing:content-box;position:absolute;top:50%;left:50%;-webkit-transform:translate(-50%,-50%);transform:translate(-50%,-50%);height:calc(100% + 4px);width:calc(100% + 4px)}@media screen and (forced-colors:active){.LQeN7 .VfPpkd-J1Ukfc-LhBDec{border-color:CanvasText}}.LQeN7 .VfPpkd-J1Ukfc-LhBDec::after{content:"";border:2px solid rgb(232,240,254);border-radius:8px;display:block;position:absolute;top:50%;left:50%;-webkit-transform:translate(-50%,-50%);transform:translate(-50%,-50%);height:calc(100% + 4px);width:calc(100% + 4px)}@media screen and (forced-colors:active){.LQeN7 .VfPpkd-J1Ukfc-LhBDec::after{border-color:CanvasText}}.LQeN7.gmghec .VfPpkd-J1Ukfc-LhBDec{display:inline-block}@media (-ms-high-contrast:active),(-ms-high-contrast:none){.LQeN7.gmghec .VfPpkd-J1Ukfc-LhBDec{display:none}}.mN1ivc .VfPpkd-Bz112c-J1Ukfc-LhBDec{pointer-events:none;border:2px solid rgb(24,90,188);border-radius:6px;box-sizing:content-box;position:absolute;top:50%;left:50%;-webkit-transform:translate(-50%,-50%);transform:translate(-50%,-50%);height:100%;width:100%}@media screen and (forced-colors:active){.mN1ivc .VfPpkd-Bz112c-J1Ukfc-LhBDec{border-color:CanvasText}}.mN1ivc .VfPpkd-Bz112c-J1Ukfc-LhBDec::after{content:"";border:2px solid rgb(232,240,254);border-radius:8px;display:block;position:absolute;top:50%;left:50%;-webkit-transform:translate(-50%,-50%);transform:translate(-50%,-50%);height:calc(100% + 4px);width:calc(100% + 4px)}@media screen and (forced-colors:active){.mN1ivc .VfPpkd-Bz112c-J1Ukfc-LhBDec::after{border-color:CanvasText}}.mN1ivc.gmghec .VfPpkd-Bz112c-J1Ukfc-LhBDec{display:inline-block}@media (-ms-high-contrast:active),(-ms-high-contrast:none){.mN1ivc.gmghec .VfPpkd-Bz112c-J1Ukfc-LhBDec{display:none}}.MyRpB .VfPpkd-kBDsod,.MyRpB .VfPpkd-vQzf8d{opacity:0}[data-tooltip-enabled=true]:disabled,.VfPpkd-Bz112c-LgbsSe[data-tooltip-enabled=true]:disabled .VfPpkd-Bz112c-Jh9lGc{pointer-events:auto}.VfPpkd-StrnGf-rymPhb{-moz-osx-font-smoothing:grayscale;-webkit-font-smoothing:antialiased;font-family:Roboto,sans-serif;font-family:var(--mdc-typography-subtitle1-font-family,var(--mdc-typography-font-family,Roboto,sans-serif));font-size:1rem;font-size:var(--mdc-typography-subtitle1-font-size,1rem);line-height:1.75rem;line-height:var(--mdc-typography-subtitle1-line-height,1.75rem);font-weight:400;font-weight:var(--mdc-typography-subtitle1-font-weight,400);letter-spacing:.009375em;letter-spacing:var(--mdc-typography-subtitle1-letter-spacing,.009375em);text-decoration:inherit;-webkit-text-decoration:var(--mdc-typography-subtitle1-text-decoration,inherit);text-decoration:var(--mdc-typography-subtitle1-text-decoration,inherit);text-transform:inherit;text-transform:var(--mdc-typography-subtitle1-text-transform,inherit);line-height:1.5rem;margin:0;padding:8px 0;list-style-type:none;color:rgba(0,0,0,.87);color:var(--mdc-theme-text-primary-on-background,rgba(0,0,0,.87))}.VfPpkd-StrnGf-rymPhb:focus{outline:none}.VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS{color:rgba(0,0,0,.54);color:var(--mdc-theme-text-secondary-on-background,rgba(0,0,0,.54))}.VfPpkd-StrnGf-rymPhb-f7MjDc{background-color:transparent}.VfPpkd-StrnGf-rymPhb-f7MjDc{color:rgba(0,0,0,.38);color:var(--mdc-theme-text-icon-on-background,rgba(0,0,0,.38))}.VfPpkd-StrnGf-rymPhb-IhFlZd{color:rgba(0,0,0,.38);color:var(--mdc-theme-text-hint-on-background,rgba(0,0,0,.38))}.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c{opacity:.38}.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS{color:#000;color:var(--mdc-theme-on-surface,#000)}.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd,.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b{color:#6200ee;color:var(--mdc-theme-primary,#6200ee)}.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-f7MjDc,.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-f7MjDc{color:#6200ee;color:var(--mdc-theme-primary,#6200ee)}.VfPpkd-StrnGf-rymPhb-OWXEXe-EzIYc{padding-top:4px;padding-bottom:4px;font-size:.812rem}.VfPpkd-StrnGf-rymPhb-Tkg0ld{display:block}.VfPpkd-StrnGf-rymPhb-Zmlebc-LhBDec{position:absolute}.VfPpkd-StrnGf-rymPhb-ibnC6b{display:-webkit-box;display:-webkit-flex;display:flex;position:relative;-webkit-box-align:center;-webkit-align-items:center;align-items:center;-webkit-box-pack:start;-webkit-justify-content:flex-start;justify-content:flex-start;overflow:hidden;padding:0;padding-left:16px;padding-right:16px;height:48px}.VfPpkd-StrnGf-rymPhb-ibnC6b:focus{outline:none}.VfPpkd-StrnGf-rymPhb-ibnC6b:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd):focus::before,.VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe::before{position:absolute;box-sizing:border-box;width:100%;height:100%;top:0;left:0;border:1px solid transparent;border-radius:inherit;content:"";pointer-events:none}@media screen and (forced-colors:active){.VfPpkd-StrnGf-rymPhb-ibnC6b:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd):focus::before,.VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe::before{border-color:CanvasText}}.VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd::before{position:absolute;box-sizing:border-box;width:100%;height:100%;top:0;left:0;border:3px double transparent;border-radius:inherit;content:"";pointer-events:none}@media screen and (forced-colors:active){.VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd::before{border-color:CanvasText}}[dir=rtl] .VfPpkd-StrnGf-rymPhb-ibnC6b,.VfPpkd-StrnGf-rymPhb-ibnC6b[dir=rtl]{padding-left:16px;padding-right:16px}.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b{padding-left:16px;padding-right:16px;height:56px}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b,.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b[dir=rtl]{padding-left:16px;padding-right:16px}.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b{padding-left:16px;padding-right:16px;height:56px}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b,.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b[dir=rtl]{padding-left:16px;padding-right:16px}.VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b{padding-left:16px;padding-right:16px;height:56px}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b,.VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b[dir=rtl]{padding-left:16px;padding-right:16px}.VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b{padding-left:16px;padding-right:16px;height:72px}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b,.VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b[dir=rtl]{padding-left:16px;padding-right:16px}.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b{padding-left:0;padding-right:16px;height:72px}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b,.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b[dir=rtl]{padding-left:16px;padding-right:0}.VfPpkd-StrnGf-rymPhb-OWXEXe-EzIYc .VfPpkd-StrnGf-rymPhb-f7MjDc{margin-left:0;margin-right:16px;width:20px;height:20px}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-EzIYc .VfPpkd-StrnGf-rymPhb-f7MjDc,.VfPpkd-StrnGf-rymPhb-OWXEXe-EzIYc .VfPpkd-StrnGf-rymPhb-f7MjDc[dir=rtl]{margin-left:16px;margin-right:0}.VfPpkd-StrnGf-rymPhb-f7MjDc{-webkit-flex-shrink:0;flex-shrink:0;-webkit-box-align:center;-webkit-align-items:center;align-items:center;-webkit-box-pack:center;-webkit-justify-content:center;justify-content:center;fill:currentColor;object-fit:cover;margin-left:0;margin-right:32px;width:24px;height:24px}[dir=rtl] .VfPpkd-StrnGf-rymPhb-f7MjDc,.VfPpkd-StrnGf-rymPhb-f7MjDc[dir=rtl]{margin-left:32px;margin-right:0}.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc{margin-left:0;margin-right:32px;width:24px;height:24px}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc,.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc[dir=rtl]{margin-left:32px;margin-right:0}.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc{margin-left:0;margin-right:16px;width:40px;height:40px;border-radius:50%}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc,.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc[dir=rtl]{margin-left:16px;margin-right:0}.VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc{margin-left:0;margin-right:16px;width:40px;height:40px}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc,.VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc[dir=rtl]{margin-left:16px;margin-right:0}.VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc{margin-left:0;margin-right:16px;width:56px;height:56px}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc,.VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc[dir=rtl]{margin-left:16px;margin-right:0}.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc{margin-left:0;margin-right:16px;width:100px;height:56px}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc,.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc[dir=rtl]{margin-left:16px;margin-right:0}.VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc{display:-webkit-inline-box;display:-webkit-inline-flex;display:inline-flex}.VfPpkd-StrnGf-rymPhb-IhFlZd{margin-left:auto;margin-right:0}.VfPpkd-StrnGf-rymPhb-IhFlZd:not(.HzV7m-fuEl3d){-moz-osx-font-smoothing:grayscale;-webkit-font-smoothing:antialiased;font-family:Roboto,sans-serif;font-family:var(--mdc-typography-caption-font-family,var(--mdc-typography-font-family,Roboto,sans-serif));font-size:.75rem;font-size:var(--mdc-typography-caption-font-size,.75rem);line-height:1.25rem;line-height:var(--mdc-typography-caption-line-height,1.25rem);font-weight:400;font-weight:var(--mdc-typography-caption-font-weight,400);letter-spacing:.0333333333em;letter-spacing:var(--mdc-typography-caption-letter-spacing,.0333333333em);text-decoration:inherit;-webkit-text-decoration:var(--mdc-typography-caption-text-decoration,inherit);text-decoration:var(--mdc-typography-caption-text-decoration,inherit);text-transform:inherit;text-transform:var(--mdc-typography-caption-text-transform,inherit)}.VfPpkd-StrnGf-rymPhb-ibnC6b[dir=rtl] .VfPpkd-StrnGf-rymPhb-IhFlZd,[dir=rtl] .VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-IhFlZd{margin-left:0;margin-right:auto}.VfPpkd-StrnGf-rymPhb-b9t22c{text-overflow:ellipsis;white-space:nowrap;overflow:hidden}.VfPpkd-StrnGf-rymPhb-b9t22c[for]{pointer-events:none}.VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS{text-overflow:ellipsis;white-space:nowrap;overflow:hidden;display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS::before{display:inline-block;width:0;height:28px;content:"";vertical-align:0}.VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS{display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS::before,.VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS::before,.VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS::before,.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS::before,.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS::before{display:inline-block;width:0;height:32px;content:"";vertical-align:0}.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS::after,.VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS::after,.VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS::after,.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS::after,.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-StrnGf-rymPhb-OWXEXe-EzIYc .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS{display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-StrnGf-rymPhb-OWXEXe-EzIYc .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS::before{display:inline-block;width:0;height:24px;content:"";vertical-align:0}.VfPpkd-StrnGf-rymPhb-OWXEXe-EzIYc .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS{-moz-osx-font-smoothing:grayscale;-webkit-font-smoothing:antialiased;font-family:Roboto,sans-serif;font-family:var(--mdc-typography-body2-font-family,var(--mdc-typography-font-family,Roboto,sans-serif));font-size:.875rem;font-size:var(--mdc-typography-body2-font-size,.875rem);line-height:1.25rem;line-height:var(--mdc-typography-body2-line-height,1.25rem);font-weight:400;font-weight:var(--mdc-typography-body2-font-weight,400);letter-spacing:.0178571429em;letter-spacing:var(--mdc-typography-body2-letter-spacing,.0178571429em);text-decoration:inherit;-webkit-text-decoration:var(--mdc-typography-body2-text-decoration,inherit);text-decoration:var(--mdc-typography-body2-text-decoration,inherit);text-transform:inherit;text-transform:var(--mdc-typography-body2-text-transform,inherit);text-overflow:ellipsis;white-space:nowrap;overflow:hidden;display:block;margin-top:0;line-height:normal}.VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS::before{display:inline-block;width:0;height:20px;content:"";vertical-align:0}.VfPpkd-StrnGf-rymPhb-OWXEXe-EzIYc .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS{font-size:inherit}.VfPpkd-StrnGf-rymPhb-OWXEXe-EzIYc .VfPpkd-StrnGf-rymPhb-ibnC6b{height:40px}.VfPpkd-StrnGf-rymPhb-OWXEXe-aSi1db-RWgCYc .VfPpkd-StrnGf-rymPhb-b9t22c{-webkit-align-self:flex-start;align-self:flex-start}.VfPpkd-StrnGf-rymPhb-OWXEXe-aSi1db-RWgCYc .VfPpkd-StrnGf-rymPhb-ibnC6b{height:64px}.VfPpkd-StrnGf-rymPhb-OWXEXe-aSi1db-RWgCYc.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b,.VfPpkd-StrnGf-rymPhb-OWXEXe-aSi1db-RWgCYc.VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b,.VfPpkd-StrnGf-rymPhb-OWXEXe-aSi1db-RWgCYc.VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b,.VfPpkd-StrnGf-rymPhb-OWXEXe-aSi1db-RWgCYc.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b,.VfPpkd-StrnGf-rymPhb-OWXEXe-aSi1db-RWgCYc.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b{height:72px}.VfPpkd-StrnGf-rymPhb-OWXEXe-aSi1db-RWgCYc.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc{-webkit-align-self:flex-start;align-self:flex-start;margin-top:16px}.VfPpkd-StrnGf-rymPhb-OWXEXe-aSi1db-RWgCYc.VfPpkd-StrnGf-rymPhb-OWXEXe-EzIYc .VfPpkd-StrnGf-rymPhb-ibnC6b,.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb.VfPpkd-StrnGf-rymPhb-OWXEXe-EzIYc .VfPpkd-StrnGf-rymPhb-ibnC6b{height:60px}.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb.VfPpkd-StrnGf-rymPhb-OWXEXe-EzIYc .VfPpkd-StrnGf-rymPhb-f7MjDc{margin-left:0;margin-right:16px;width:36px;height:36px}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb.VfPpkd-StrnGf-rymPhb-OWXEXe-EzIYc .VfPpkd-StrnGf-rymPhb-f7MjDc,.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb.VfPpkd-StrnGf-rymPhb-OWXEXe-EzIYc .VfPpkd-StrnGf-rymPhb-f7MjDc[dir=rtl]{margin-left:16px;margin-right:0}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b{cursor:pointer}a.VfPpkd-StrnGf-rymPhb-ibnC6b{color:inherit;text-decoration:none}.VfPpkd-StrnGf-rymPhb-clz4Ic{height:0;margin:0;border:none;border-bottom-width:1px;border-bottom-style:solid}.VfPpkd-StrnGf-rymPhb-clz4Ic{border-bottom-color:rgba(0,0,0,.12)}.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-nNtqDd{margin-left:16px;margin-right:0;width:calc(100% - 32px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-nNtqDd,.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-nNtqDd[dir=rtl]{margin-left:0;margin-right:16px}.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe{margin-left:72px;margin-right:0;width:calc(100% - 72px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe,.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe[dir=rtl]{margin-left:0;margin-right:72px}.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-nNtqDd{margin-left:72px;margin-right:0;width:calc(100% - 88px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-nNtqDd,.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-nNtqDd[dir=rtl]{margin-left:0;margin-right:72px}.VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc{margin-left:16px;margin-right:0;width:calc(100% - 16px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc,.VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc[dir=rtl]{margin-left:0;margin-right:16px}.VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg{width:calc(100% - 16px)}.VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg{margin-left:16px;margin-right:0;width:calc(100% - 32px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg,.VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg[dir=rtl]{margin-left:0;margin-right:16px}.VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2{margin-left:16px;margin-right:0;width:calc(100% - 16px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2,.VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2[dir=rtl]{margin-left:0;margin-right:16px}.VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2{margin-left:16px;margin-right:0;width:calc(100% - 32px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2,.VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2[dir=rtl]{margin-left:0;margin-right:16px}.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc{margin-left:72px;margin-right:0;width:calc(100% - 72px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc,.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc[dir=rtl]{margin-left:0;margin-right:72px}.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg{width:calc(100% - 16px)}.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg{margin-left:72px;margin-right:0;width:calc(100% - 88px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg,.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg[dir=rtl]{margin-left:0;margin-right:72px}.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2{margin-left:16px;margin-right:0;width:calc(100% - 16px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2,.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2[dir=rtl]{margin-left:0;margin-right:16px}.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2{margin-left:16px;margin-right:0;width:calc(100% - 32px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2,.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2[dir=rtl]{margin-left:0;margin-right:16px}.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc{margin-left:72px;margin-right:0;width:calc(100% - 72px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc,.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc[dir=rtl]{margin-left:0;margin-right:72px}.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg{width:calc(100% - 16px)}.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg{margin-left:72px;margin-right:0;width:calc(100% - 88px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg,.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg[dir=rtl]{margin-left:0;margin-right:72px}.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2{margin-left:16px;margin-right:0;width:calc(100% - 16px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2,.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2[dir=rtl]{margin-left:0;margin-right:16px}.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2{margin-left:16px;margin-right:0;width:calc(100% - 32px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2,.VfPpkd-StrnGf-rymPhb-OWXEXe-YLEF4c-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2[dir=rtl]{margin-left:0;margin-right:16px}.VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc{margin-left:72px;margin-right:0;width:calc(100% - 72px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc,.VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc[dir=rtl]{margin-left:0;margin-right:72px}.VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg{width:calc(100% - 16px)}.VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg{margin-left:72px;margin-right:0;width:calc(100% - 88px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg,.VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg[dir=rtl]{margin-left:0;margin-right:72px}.VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2{margin-left:16px;margin-right:0;width:calc(100% - 16px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2,.VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2[dir=rtl]{margin-left:0;margin-right:16px}.VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2{margin-left:16px;margin-right:0;width:calc(100% - 32px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2,.VfPpkd-StrnGf-rymPhb-OWXEXe-JUCs7e-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2[dir=rtl]{margin-left:0;margin-right:16px}.VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc{margin-left:88px;margin-right:0;width:calc(100% - 88px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc,.VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc[dir=rtl]{margin-left:0;margin-right:88px}.VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg{width:calc(100% - 16px)}.VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg{margin-left:88px;margin-right:0;width:calc(100% - 104px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg,.VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg[dir=rtl]{margin-left:0;margin-right:88px}.VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2{margin-left:16px;margin-right:0;width:calc(100% - 16px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2,.VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2[dir=rtl]{margin-left:0;margin-right:16px}.VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2{margin-left:16px;margin-right:0;width:calc(100% - 32px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2,.VfPpkd-StrnGf-rymPhb-OWXEXe-HiaYvf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2[dir=rtl]{margin-left:0;margin-right:16px}.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc{margin-left:116px;margin-right:0;width:calc(100% - 116px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc,.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc[dir=rtl]{margin-left:0;margin-right:116px}.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg{width:calc(100% - 16px)}.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg{margin-left:116px;margin-right:0;width:calc(100% - 132px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg,.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg[dir=rtl]{margin-left:0;margin-right:116px}.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2{margin-left:0;margin-right:0;width:100%}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2,.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2[dir=rtl]{margin-left:0;margin-right:0}.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2{margin-left:0;margin-right:0;width:calc(100% - 16px)}[dir=rtl] .VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2,.VfPpkd-StrnGf-rymPhb-OWXEXe-aTv5jf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2[dir=rtl]{margin-left:0;margin-right:0}.VfPpkd-StrnGf-rymPhb-JNdkSc .VfPpkd-StrnGf-rymPhb{padding:0}.VfPpkd-StrnGf-rymPhb-oT7voc{-moz-osx-font-smoothing:grayscale;-webkit-font-smoothing:antialiased;font-family:Roboto,sans-serif;font-family:var(--mdc-typography-subtitle1-font-family,var(--mdc-typography-font-family,Roboto,sans-serif));font-size:1rem;font-size:var(--mdc-typography-subtitle1-font-size,1rem);line-height:1.75rem;line-height:var(--mdc-typography-subtitle1-line-height,1.75rem);font-weight:400;font-weight:var(--mdc-typography-subtitle1-font-weight,400);letter-spacing:.009375em;letter-spacing:var(--mdc-typography-subtitle1-letter-spacing,.009375em);text-decoration:inherit;-webkit-text-decoration:var(--mdc-typography-subtitle1-text-decoration,inherit);text-decoration:var(--mdc-typography-subtitle1-text-decoration,inherit);text-transform:inherit;text-transform:var(--mdc-typography-subtitle1-text-transform,inherit);margin:.75rem 16px}.VfPpkd-rymPhb-Gtdoyb,.VfPpkd-rymPhb-fpDzbe-fmcmS{color:rgba(0,0,0,.87);color:var(--mdc-theme-text-primary-on-background,rgba(0,0,0,.87))}.VfPpkd-rymPhb-L8ivfd-fmcmS{color:rgba(0,0,0,.54);color:var(--mdc-theme-text-secondary-on-background,rgba(0,0,0,.54))}.VfPpkd-rymPhb-bC5pod-fmcmS{color:rgba(0,0,0,.38);color:var(--mdc-theme-text-hint-on-background,rgba(0,0,0,.38))}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e{background-color:transparent}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e{color:rgba(0,0,0,.38);color:var(--mdc-theme-text-icon-on-background,rgba(0,0,0,.38))}.VfPpkd-rymPhb-JMEf7e{color:rgba(0,0,0,.38);color:var(--mdc-theme-text-hint-on-background,rgba(0,0,0,.38))}.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-KkROqb,.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-Gtdoyb,.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-JMEf7e{opacity:.38}.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-Gtdoyb,.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-fpDzbe-fmcmS{color:#000;color:var(--mdc-theme-on-surface,#000)}.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-L8ivfd-fmcmS{color:#000;color:var(--mdc-theme-on-surface,#000)}.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-bC5pod-fmcmS{color:#000;color:var(--mdc-theme-on-surface,#000)}.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb{color:#000;color:var(--mdc-theme-on-surface,#000)}.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e{color:#000;color:var(--mdc-theme-on-surface,#000)}.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e{color:#000;color:var(--mdc-theme-on-surface,#000)}.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-Gtdoyb,.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-fpDzbe-fmcmS,.VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-rymPhb-Gtdoyb,.VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-rymPhb-fpDzbe-fmcmS{color:#6200ee;color:var(--mdc-theme-primary,#6200ee)}.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb,.VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb{color:#6200ee;color:var(--mdc-theme-primary,#6200ee)}.VfPpkd-StrnGf-rymPhb-oT7voc{color:rgba(0,0,0,.87);color:var(--mdc-theme-text-primary-on-background,rgba(0,0,0,.87))}.VfPpkd-rymPhb-clz4Ic::after{border-bottom-color:white}.VfPpkd-rymPhb{-moz-osx-font-smoothing:grayscale;-webkit-font-smoothing:antialiased;font-family:Roboto,sans-serif;font-family:var(--mdc-typography-subtitle1-font-family,var(--mdc-typography-font-family,Roboto,sans-serif));font-size:1rem;font-size:var(--mdc-typography-subtitle1-font-size,1rem);line-height:1.75rem;line-height:var(--mdc-typography-subtitle1-line-height,1.75rem);font-weight:400;font-weight:var(--mdc-typography-subtitle1-font-weight,400);letter-spacing:.009375em;letter-spacing:var(--mdc-typography-subtitle1-letter-spacing,.009375em);text-decoration:inherit;-webkit-text-decoration:var(--mdc-typography-subtitle1-text-decoration,inherit);text-decoration:var(--mdc-typography-subtitle1-text-decoration,inherit);text-transform:inherit;text-transform:var(--mdc-typography-subtitle1-text-transform,inherit);line-height:1.5rem}.VfPpkd-rymPhb-fpDzbe-fmcmS{-moz-osx-font-smoothing:grayscale;-webkit-font-smoothing:antialiased;font-family:Roboto,sans-serif;font-family:var(--mdc-typography-subtitle1-font-family,var(--mdc-typography-font-family,Roboto,sans-serif));font-size:1rem;font-size:var(--mdc-typography-subtitle1-font-size,1rem);line-height:1.75rem;line-height:var(--mdc-typography-subtitle1-line-height,1.75rem);font-weight:400;font-weight:var(--mdc-typography-subtitle1-font-weight,400);letter-spacing:.009375em;letter-spacing:var(--mdc-typography-subtitle1-letter-spacing,.009375em);text-decoration:inherit;-webkit-text-decoration:var(--mdc-typography-subtitle1-text-decoration,inherit);text-decoration:var(--mdc-typography-subtitle1-text-decoration,inherit);text-transform:inherit;text-transform:var(--mdc-typography-subtitle1-text-transform,inherit)}.VfPpkd-rymPhb-L8ivfd-fmcmS{-moz-osx-font-smoothing:grayscale;-webkit-font-smoothing:antialiased;font-family:Roboto,sans-serif;font-family:var(--mdc-typography-body2-font-family,var(--mdc-typography-font-family,Roboto,sans-serif));font-size:.875rem;font-size:var(--mdc-typography-body2-font-size,.875rem);line-height:1.25rem;line-height:var(--mdc-typography-body2-line-height,1.25rem);font-weight:400;font-weight:var(--mdc-typography-body2-font-weight,400);letter-spacing:.0178571429em;letter-spacing:var(--mdc-typography-body2-letter-spacing,.0178571429em);text-decoration:inherit;-webkit-text-decoration:var(--mdc-typography-body2-text-decoration,inherit);text-decoration:var(--mdc-typography-body2-text-decoration,inherit);text-transform:inherit;text-transform:var(--mdc-typography-body2-text-transform,inherit)}.VfPpkd-rymPhb-bC5pod-fmcmS{-moz-osx-font-smoothing:grayscale;-webkit-font-smoothing:antialiased;font-family:Roboto,sans-serif;font-family:var(--mdc-typography-overline-font-family,var(--mdc-typography-font-family,Roboto,sans-serif));font-size:.75rem;font-size:var(--mdc-typography-overline-font-size,.75rem);line-height:2rem;line-height:var(--mdc-typography-overline-line-height,2rem);font-weight:500;font-weight:var(--mdc-typography-overline-font-weight,500);letter-spacing:.1666666667em;letter-spacing:var(--mdc-typography-overline-letter-spacing,.1666666667em);text-decoration:none;-webkit-text-decoration:var(--mdc-typography-overline-text-decoration,none);text-decoration:var(--mdc-typography-overline-text-decoration,none);text-transform:uppercase;text-transform:var(--mdc-typography-overline-text-transform,uppercase)}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c .VfPpkd-rymPhb-KkROqb{width:40px;height:40px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb{width:24px;height:24px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e .VfPpkd-rymPhb-KkROqb{width:40px;height:40px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf .VfPpkd-rymPhb-KkROqb{width:56px;height:56px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf .VfPpkd-rymPhb-KkROqb{width:100px;height:56px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c .VfPpkd-rymPhb-KkROqb,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b .VfPpkd-rymPhb-KkROqb{width:40px;height:40px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc .VfPpkd-rymPhb-KkROqb{width:36px;height:20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e{width:24px;height:24px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-MPu53c .VfPpkd-rymPhb-JMEf7e,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-GCYh9b .VfPpkd-rymPhb-JMEf7e{width:40px;height:40px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-scr2fc .VfPpkd-rymPhb-JMEf7e{width:36px;height:20px}.VfPpkd-rymPhb-oT7voc{-moz-osx-font-smoothing:grayscale;-webkit-font-smoothing:antialiased;font-family:Roboto,sans-serif;font-family:var(--mdc-typography-subtitle1-font-family,var(--mdc-typography-font-family,Roboto,sans-serif));font-size:1rem;font-size:var(--mdc-typography-subtitle1-font-size,1rem);line-height:1.75rem;line-height:var(--mdc-typography-subtitle1-line-height,1.75rem);font-weight:400;font-weight:var(--mdc-typography-subtitle1-font-weight,400);letter-spacing:.009375em;letter-spacing:var(--mdc-typography-subtitle1-letter-spacing,.009375em);text-decoration:inherit;-webkit-text-decoration:var(--mdc-typography-subtitle1-text-decoration,inherit);text-decoration:var(--mdc-typography-subtitle1-text-decoration,inherit);text-transform:inherit;text-transform:var(--mdc-typography-subtitle1-text-transform,inherit)}.VfPpkd-rymPhb-clz4Ic{background-color:rgba(0,0,0,.12)}.VfPpkd-rymPhb-clz4Ic{height:1px}@media (-ms-high-contrast:active),screen and (forced-colors:active){.VfPpkd-rymPhb-clz4Ic::after{content:"";display:block;border-bottom-width:1px;border-bottom-style:solid}}.VfPpkd-rymPhb{margin:0;padding:8px 0;list-style-type:none}.VfPpkd-rymPhb:focus{outline:none}.VfPpkd-rymPhb-Tkg0ld{display:block}.VfPpkd-rymPhb-ibnC6b{display:-webkit-box;display:-webkit-flex;display:flex;position:relative;-webkit-box-align:center;-webkit-align-items:center;align-items:center;-webkit-box-pack:start;-webkit-justify-content:flex-start;justify-content:flex-start;overflow:hidden;padding:0;-webkit-box-align:stretch;-webkit-align-items:stretch;align-items:stretch;cursor:pointer}.VfPpkd-rymPhb-ibnC6b:focus{outline:none}.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc{height:48px}.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb{height:64px}.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb{height:88px}.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc .VfPpkd-rymPhb-KkROqb{-webkit-align-self:center;align-self:center;margin-top:0}.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-KkROqb,.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-KkROqb{-webkit-align-self:flex-start;align-self:flex-start;margin-top:16px}.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc .VfPpkd-rymPhb-JMEf7e,.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-JMEf7e{-webkit-align-self:center;align-self:center;margin-top:0}.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-JMEf7e{-webkit-align-self:flex-start;align-self:flex-start;margin-top:16px}.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me,.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-tPcied-hXIJHe{cursor:auto}.VfPpkd-rymPhb-ibnC6b:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd):focus::before,.VfPpkd-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe::before{position:absolute;box-sizing:border-box;width:100%;height:100%;top:0;left:0;border:1px solid transparent;border-radius:inherit;content:"";pointer-events:none}@media screen and (forced-colors:active){.VfPpkd-rymPhb-ibnC6b:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd):focus::before,.VfPpkd-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe::before{border-color:CanvasText}}.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd::before{position:absolute;box-sizing:border-box;width:100%;height:100%;top:0;left:0;border:3px double transparent;border-radius:inherit;content:"";pointer-events:none}@media screen and (forced-colors:active){.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd::before{border-color:CanvasText}}.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:focus::before{position:absolute;box-sizing:border-box;width:100%;height:100%;top:0;left:0;border:3px solid transparent;border-radius:inherit;content:"";pointer-events:none}@media screen and (forced-colors:active){.VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:focus::before{border-color:CanvasText}}a.VfPpkd-rymPhb-ibnC6b{color:inherit;text-decoration:none}.VfPpkd-rymPhb-KkROqb{fill:currentColor;-webkit-flex-shrink:0;flex-shrink:0;pointer-events:none}.VfPpkd-rymPhb-JMEf7e{-webkit-flex-shrink:0;flex-shrink:0;pointer-events:none}.VfPpkd-rymPhb-Gtdoyb{text-overflow:ellipsis;white-space:nowrap;overflow:hidden;-webkit-align-self:center;align-self:center;-webkit-box-flex:1;-webkit-flex:1;flex:1;pointer-events:none}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-Gtdoyb,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-Gtdoyb{-webkit-align-self:stretch;align-self:stretch}.VfPpkd-rymPhb-Gtdoyb[for]{pointer-events:none}.VfPpkd-rymPhb-fpDzbe-fmcmS{text-overflow:ellipsis;white-space:nowrap;overflow:hidden}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS{display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::before,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::before{display:inline-block;width:0;height:28px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::after,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-rymPhb-L8ivfd-fmcmS{text-overflow:ellipsis;white-space:nowrap;overflow:hidden;display:block;margin-top:0;line-height:normal}.VfPpkd-rymPhb-L8ivfd-fmcmS::before{display:inline-block;width:0;height:20px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-L8ivfd-fmcmS{white-space:normal;line-height:20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-BYmFj .VfPpkd-rymPhb-L8ivfd-fmcmS{white-space:nowrap;line-height:auto}.VfPpkd-rymPhb-bC5pod-fmcmS{text-overflow:ellipsis;white-space:nowrap;overflow:hidden}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS{display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::before{display:inline-block;width:0;height:24px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS{display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::before{display:inline-block;width:0;height:28px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-ibnC6b{padding-left:0;padding-right:auto}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-ibnC6b,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:auto;padding-right:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c .VfPpkd-rymPhb-KkROqb{margin-left:16px;margin-right:16px}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c .VfPpkd-rymPhb-KkROqb,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c .VfPpkd-rymPhb-KkROqb[dir=rtl]{margin-left:16px;margin-right:16px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS{display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::before{display:inline-block;width:0;height:32px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS{display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::before{display:inline-block;width:0;height:28px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e{display:block;margin-top:0;line-height:normal}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e::before{display:inline-block;width:0;height:32px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc{height:56px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb{height:72px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-YLEF4c .VfPpkd-rymPhb-KkROqb{border-radius:50%}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-ibnC6b{padding-left:0;padding-right:auto}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-ibnC6b,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:auto;padding-right:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb{margin-left:16px;margin-right:32px}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb[dir=rtl]{margin-left:32px;margin-right:16px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS{display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::before{display:inline-block;width:0;height:32px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS{display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::before{display:inline-block;width:0;height:28px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e{display:block;margin-top:0;line-height:normal}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e::before{display:inline-block;width:0;height:32px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc{height:56px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb{height:72px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-ibnC6b{padding-left:0;padding-right:auto}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-ibnC6b,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:auto;padding-right:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e .VfPpkd-rymPhb-KkROqb{margin-left:16px;margin-right:16px}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e .VfPpkd-rymPhb-KkROqb,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e .VfPpkd-rymPhb-KkROqb[dir=rtl]{margin-left:16px;margin-right:16px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS{display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::before{display:inline-block;width:0;height:32px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS{display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::before{display:inline-block;width:0;height:28px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e{display:block;margin-top:0;line-height:normal}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e::before{display:inline-block;width:0;height:32px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc{height:56px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb{height:72px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b{padding-left:0;padding-right:auto}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:auto;padding-right:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf .VfPpkd-rymPhb-KkROqb{margin-left:16px;margin-right:16px}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf .VfPpkd-rymPhb-KkROqb,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf .VfPpkd-rymPhb-KkROqb[dir=rtl]{margin-left:16px;margin-right:16px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS{display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::before{display:inline-block;width:0;height:32px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS{display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::before{display:inline-block;width:0;height:28px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e{display:block;margin-top:0;line-height:normal}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e::before{display:inline-block;width:0;height:32px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb{height:72px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-KkROqb{-webkit-align-self:flex-start;align-self:flex-start;margin-top:8px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b{padding-left:0;padding-right:auto}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:auto;padding-right:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf .VfPpkd-rymPhb-KkROqb{margin-left:0;margin-right:16px}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf .VfPpkd-rymPhb-KkROqb,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf .VfPpkd-rymPhb-KkROqb[dir=rtl]{margin-left:16px;margin-right:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS{display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::before{display:inline-block;width:0;height:32px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS{display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::before{display:inline-block;width:0;height:28px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e{display:block;margin-top:0;line-height:normal}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e::before{display:inline-block;width:0;height:32px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb{height:72px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b{padding-left:0;padding-right:auto}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:auto;padding-right:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c .VfPpkd-rymPhb-KkROqb{margin-left:8px;margin-right:24px}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c .VfPpkd-rymPhb-KkROqb,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c .VfPpkd-rymPhb-KkROqb[dir=rtl]{margin-left:24px;margin-right:8px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-KkROqb{-webkit-align-self:flex-start;align-self:flex-start;margin-top:8px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS{display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::before{display:inline-block;width:0;height:32px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS{display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::before{display:inline-block;width:0;height:28px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e{display:block;margin-top:0;line-height:normal}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e::before{display:inline-block;width:0;height:32px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc{height:56px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb{height:72px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b{padding-left:0;padding-right:auto}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:auto;padding-right:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b .VfPpkd-rymPhb-KkROqb{margin-left:8px;margin-right:24px}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b .VfPpkd-rymPhb-KkROqb,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b .VfPpkd-rymPhb-KkROqb[dir=rtl]{margin-left:24px;margin-right:8px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-KkROqb{-webkit-align-self:flex-start;align-self:flex-start;margin-top:8px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS{display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::before{display:inline-block;width:0;height:32px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS{display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::before{display:inline-block;width:0;height:28px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e{display:block;margin-top:0;line-height:normal}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e::before{display:inline-block;width:0;height:32px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc{height:56px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb{height:72px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b{padding-left:0;padding-right:auto}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:auto;padding-right:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc .VfPpkd-rymPhb-KkROqb{margin-left:16px;margin-right:16px}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc .VfPpkd-rymPhb-KkROqb,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc .VfPpkd-rymPhb-KkROqb[dir=rtl]{margin-left:16px;margin-right:16px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-KkROqb{-webkit-align-self:flex-start;align-self:flex-start;margin-top:16px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS{display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::before{display:inline-block;width:0;height:32px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS{display:block;margin-top:0;line-height:normal;margin-bottom:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::before{display:inline-block;width:0;height:28px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-bC5pod-fmcmS::after{display:inline-block;width:0;height:20px;content:"";vertical-align:-20px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e{display:block;margin-top:0;line-height:normal}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e::before{display:inline-block;width:0;height:32px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc{height:56px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb{height:72px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c.VfPpkd-rymPhb-ibnC6b{padding-left:auto;padding-right:0}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c.VfPpkd-rymPhb-ibnC6b,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:0;padding-right:auto}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e{margin-left:16px;margin-right:16px}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e[dir=rtl]{margin-left:16px;margin-right:16px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-JMEf7e,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-JMEf7e{-webkit-align-self:flex-start;align-self:flex-start;margin-top:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf.VfPpkd-rymPhb-ibnC6b{padding-left:auto;padding-right:0}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf.VfPpkd-rymPhb-ibnC6b,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:0;padding-right:auto}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e{margin-left:28px;margin-right:16px}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e[dir=rtl]{margin-left:16px;margin-right:28px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-JMEf7e{display:block;margin-top:0;line-height:normal}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-JMEf7e::before{display:inline-block;width:0;height:28px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-JMEf7e{display:block;margin-top:0;line-height:normal}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-JMEf7e::before{display:inline-block;width:0;height:28px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e{-moz-osx-font-smoothing:grayscale;-webkit-font-smoothing:antialiased;font-family:Roboto,sans-serif;font-family:var(--mdc-typography-caption-font-family,var(--mdc-typography-font-family,Roboto,sans-serif));font-size:.75rem;font-size:var(--mdc-typography-caption-font-size,.75rem);line-height:1.25rem;line-height:var(--mdc-typography-caption-line-height,1.25rem);font-weight:400;font-weight:var(--mdc-typography-caption-font-weight,400);letter-spacing:.0333333333em;letter-spacing:var(--mdc-typography-caption-letter-spacing,.0333333333em);text-decoration:inherit;-webkit-text-decoration:var(--mdc-typography-caption-text-decoration,inherit);text-decoration:var(--mdc-typography-caption-text-decoration,inherit);text-transform:inherit;text-transform:var(--mdc-typography-caption-text-transform,inherit)}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-MPu53c.VfPpkd-rymPhb-ibnC6b{padding-left:auto;padding-right:0}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-MPu53c.VfPpkd-rymPhb-ibnC6b,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-MPu53c.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:0;padding-right:auto}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-MPu53c .VfPpkd-rymPhb-JMEf7e{margin-left:24px;margin-right:8px}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-MPu53c .VfPpkd-rymPhb-JMEf7e,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-MPu53c .VfPpkd-rymPhb-JMEf7e[dir=rtl]{margin-left:8px;margin-right:24px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-MPu53c.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-JMEf7e{-webkit-align-self:flex-start;align-self:flex-start;margin-top:8px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-GCYh9b.VfPpkd-rymPhb-ibnC6b{padding-left:auto;padding-right:0}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-GCYh9b.VfPpkd-rymPhb-ibnC6b,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-GCYh9b.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:0;padding-right:auto}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-GCYh9b .VfPpkd-rymPhb-JMEf7e{margin-left:24px;margin-right:8px}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-GCYh9b .VfPpkd-rymPhb-JMEf7e,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-GCYh9b .VfPpkd-rymPhb-JMEf7e[dir=rtl]{margin-left:8px;margin-right:24px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-GCYh9b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-JMEf7e{-webkit-align-self:flex-start;align-self:flex-start;margin-top:8px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-scr2fc.VfPpkd-rymPhb-ibnC6b{padding-left:auto;padding-right:0}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-scr2fc.VfPpkd-rymPhb-ibnC6b,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-scr2fc.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:0;padding-right:auto}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-scr2fc .VfPpkd-rymPhb-JMEf7e{margin-left:16px;margin-right:16px}[dir=rtl] .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-scr2fc .VfPpkd-rymPhb-JMEf7e,.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-scr2fc .VfPpkd-rymPhb-JMEf7e[dir=rtl]{margin-left:16px;margin-right:16px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-scr2fc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-JMEf7e{-webkit-align-self:flex-start;align-self:flex-start;margin-top:16px}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-BYmFj.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS{display:block;margin-top:0;line-height:normal}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-BYmFj.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::before{display:inline-block;width:0;height:20px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-BYmFj.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS{display:block;margin-top:0;line-height:normal}.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-BYmFj.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-vfifzc-MCEKJb .VfPpkd-rymPhb-fpDzbe-fmcmS::before{display:inline-block;width:0;height:20px;content:"";vertical-align:0}.VfPpkd-rymPhb-ibnC6b{padding-left:16px;padding-right:16px}[dir=rtl] .VfPpkd-rymPhb-ibnC6b,.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:16px;padding-right:16px}.VfPpkd-rymPhb-JNdkSc .VfPpkd-StrnGf-rymPhb{padding:0}.VfPpkd-rymPhb-oT7voc{margin:.75rem 16px}.VfPpkd-rymPhb-clz4Ic{padding:0;background-clip:content-box}.VfPpkd-rymPhb-clz4Ic.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe,.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-fmcmS.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe,.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe,.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe,.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe,.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe,.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe,.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe,.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe{padding-left:16px;padding-right:auto}[dir=rtl] .VfPpkd-rymPhb-clz4Ic.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe,[dir=rtl] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-fmcmS.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe,[dir=rtl] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe,[dir=rtl] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe,[dir=rtl] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe,[dir=rtl] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe,[dir=rtl] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe,[dir=rtl] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe,[dir=rtl] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe,.VfPpkd-rymPhb-clz4Ic.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe[dir=rtl],.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-fmcmS.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe[dir=rtl],.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe[dir=rtl],.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe[dir=rtl],.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe[dir=rtl],.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe[dir=rtl],.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe[dir=rtl],.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe[dir=rtl],.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe[dir=rtl]{padding-left:auto;padding-right:16px}.VfPpkd-rymPhb-clz4Ic.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe,.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-fmcmS.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe,.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe,.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe,.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe,.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe,.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe,.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe,.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe{padding-left:auto;padding-right:16px}[dir=rtl] .VfPpkd-rymPhb-clz4Ic.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe,[dir=rtl] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-fmcmS.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe,[dir=rtl] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe,[dir=rtl] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe,[dir=rtl] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe,[dir=rtl] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe,[dir=rtl] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe,[dir=rtl] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe,[dir=rtl] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe,.VfPpkd-rymPhb-clz4Ic.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe[dir=rtl],.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-fmcmS.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe[dir=rtl],.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-Bz112c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe[dir=rtl],.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe[dir=rtl],.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-JUCs7e.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe[dir=rtl],.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YLEF4c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe[dir=rtl],.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-MPu53c.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe[dir=rtl],.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-scr2fc.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe[dir=rtl],.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-GCYh9b.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe[dir=rtl]{padding-left:16px;padding-right:auto}.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe{padding-left:0;padding-right:auto}[dir=rtl] .VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe,.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe[dir=rtl]{padding-left:auto;padding-right:0}[dir=rtl] .VfPpkd-rymPhb-clz4Ic,.VfPpkd-rymPhb-clz4Ic[dir=rtl]{padding:0}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b{--mdc-ripple-fg-size:0;--mdc-ripple-left:0;--mdc-ripple-top:0;--mdc-ripple-fg-scale:1;--mdc-ripple-fg-translate-end:0;--mdc-ripple-fg-translate-start:0;-webkit-tap-highlight-color:rgba(0,0,0,0);will-change:transform,opacity}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-pZXsl::before,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-pZXsl::after{position:absolute;border-radius:50%;opacity:0;pointer-events:none;content:""}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-pZXsl::before{-webkit-transition:opacity 15ms linear,background-color 15ms linear;transition:opacity 15ms linear,background-color 15ms linear;z-index:1;z-index:var(--mdc-ripple-z-index,1)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-pZXsl::after{z-index:0;z-index:var(--mdc-ripple-z-index,0)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d .VfPpkd-StrnGf-rymPhb-pZXsl::before{-webkit-transform:scale(var(--mdc-ripple-fg-scale,1));transform:scale(var(--mdc-ripple-fg-scale,1))}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d .VfPpkd-StrnGf-rymPhb-pZXsl::after{top:0;left:0;-webkit-transform:scale(0);transform:scale(0);-webkit-transform-origin:center center;transform-origin:center center}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd .VfPpkd-StrnGf-rymPhb-pZXsl::after{top:var(--mdc-ripple-top,0);left:var(--mdc-ripple-left,0)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-lJfZMc .VfPpkd-StrnGf-rymPhb-pZXsl::after{-webkit-animation:mdc-ripple-fg-radius-in 225ms forwards,mdc-ripple-fg-opacity-in 75ms forwards;animation:mdc-ripple-fg-radius-in 225ms forwards,mdc-ripple-fg-opacity-in 75ms forwards}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-OmS1vf .VfPpkd-StrnGf-rymPhb-pZXsl::after{-webkit-animation:mdc-ripple-fg-opacity-out .15s;animation:mdc-ripple-fg-opacity-out .15s;-webkit-transform:translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1));transform:translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1))}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::before,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::after{position:absolute;border-radius:50%;opacity:0;pointer-events:none;content:""}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::before{-webkit-transition:opacity 15ms linear,background-color 15ms linear;transition:opacity 15ms linear,background-color 15ms linear;z-index:1;z-index:var(--mdc-ripple-z-index,1)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::after{z-index:0;z-index:var(--mdc-ripple-z-index,0)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d .VfPpkd-rymPhb-pZXsl::before{-webkit-transform:scale(var(--mdc-ripple-fg-scale,1));transform:scale(var(--mdc-ripple-fg-scale,1))}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d .VfPpkd-rymPhb-pZXsl::after{top:0;left:0;-webkit-transform:scale(0);transform:scale(0);-webkit-transform-origin:center center;transform-origin:center center}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd .VfPpkd-rymPhb-pZXsl::after{top:var(--mdc-ripple-top,0);left:var(--mdc-ripple-left,0)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-lJfZMc .VfPpkd-rymPhb-pZXsl::after{-webkit-animation:mdc-ripple-fg-radius-in 225ms forwards,mdc-ripple-fg-opacity-in 75ms forwards;animation:mdc-ripple-fg-radius-in 225ms forwards,mdc-ripple-fg-opacity-in 75ms forwards}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-OmS1vf .VfPpkd-rymPhb-pZXsl::after{-webkit-animation:mdc-ripple-fg-opacity-out .15s;animation:mdc-ripple-fg-opacity-out .15s;-webkit-transform:translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1));transform:translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1))}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-pZXsl::before,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-pZXsl::after{top:-50%;left:-50%;width:200%;height:200%}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d .VfPpkd-StrnGf-rymPhb-pZXsl::after{width:var(--mdc-ripple-fg-size,100%);height:var(--mdc-ripple-fg-size,100%)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::before,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::after{top:-50%;left:-50%;width:200%;height:200%}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d .VfPpkd-rymPhb-pZXsl::after{width:var(--mdc-ripple-fg-size,100%);height:var(--mdc-ripple-fg-size,100%)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-pZXsl::before,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-pZXsl::after{background-color:#000;background-color:var(--mdc-ripple-color,#000)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-press-opacity,.12)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::before,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::after{background-color:#000;background-color:var(--mdc-ripple-color,#000)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b:hover .VfPpkd-rymPhb-pZXsl::before,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-rymPhb-pZXsl::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-rymPhb-pZXsl::before,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-rymPhb-pZXsl::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-rymPhb-pZXsl::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-rymPhb-pZXsl::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-press-opacity,.12)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.12)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:.12;opacity:var(--mdc-ripple-activated-opacity,.12)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-pZXsl::before,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-pZXsl::after{background-color:#6200ee;background-color:var(--mdc-ripple-color,var(--mdc-theme-primary,#6200ee))}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:.16;opacity:var(--mdc-ripple-hover-opacity,.16)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.24;opacity:var(--mdc-ripple-focus-opacity,.24)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.24;opacity:var(--mdc-ripple-press-opacity,.24)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-rymPhb-pZXsl::before{opacity:.12;opacity:var(--mdc-ripple-activated-opacity,.12)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-rymPhb-pZXsl::before,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-rymPhb-pZXsl::after{background-color:#6200ee;background-color:var(--mdc-ripple-color,var(--mdc-theme-primary,#6200ee))}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b:hover .VfPpkd-rymPhb-pZXsl::before,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-rymPhb-pZXsl::before{opacity:.16;opacity:var(--mdc-ripple-hover-opacity,.16)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-rymPhb-pZXsl::before,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-rymPhb-pZXsl::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.24;opacity:var(--mdc-ripple-focus-opacity,.24)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-rymPhb-pZXsl::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-rymPhb-pZXsl::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.24;opacity:var(--mdc-ripple-press-opacity,.24)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.24)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:.08;opacity:var(--mdc-ripple-selected-opacity,.08)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::after{background-color:#6200ee;background-color:var(--mdc-ripple-color,var(--mdc-theme-primary,#6200ee))}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:.12;opacity:var(--mdc-ripple-hover-opacity,.12)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.2;opacity:var(--mdc-ripple-focus-opacity,.2)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.2;opacity:var(--mdc-ripple-press-opacity,.2)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::before{opacity:.08;opacity:var(--mdc-ripple-selected-opacity,.08)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::before,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::after{background-color:#6200ee;background-color:var(--mdc-ripple-color,var(--mdc-theme-primary,#6200ee))}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-rymPhb-pZXsl::before,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-rymPhb-pZXsl::before{opacity:.12;opacity:var(--mdc-ripple-hover-opacity,.12)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-rymPhb-pZXsl::before,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-rymPhb-pZXsl::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.2;opacity:var(--mdc-ripple-focus-opacity,.2)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-rymPhb-pZXsl::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-rymPhb-pZXsl::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.2;opacity:var(--mdc-ripple-press-opacity,.2)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.2)}:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-pZXsl,:not(.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl{position:absolute;top:0;left:0;width:100%;height:100%;pointer-events:none}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b{--mdc-ripple-fg-size:0;--mdc-ripple-left:0;--mdc-ripple-top:0;--mdc-ripple-fg-scale:1;--mdc-ripple-fg-translate-end:0;--mdc-ripple-fg-translate-start:0;-webkit-tap-highlight-color:rgba(0,0,0,0);will-change:transform,opacity}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::before,:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::after{position:absolute;border-radius:50%;opacity:0;pointer-events:none;content:""}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::before{-webkit-transition:opacity 15ms linear,background-color 15ms linear;transition:opacity 15ms linear,background-color 15ms linear;z-index:1;z-index:var(--mdc-ripple-z-index,1)}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::after{z-index:0;z-index:var(--mdc-ripple-z-index,0)}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d .VfPpkd-rymPhb-pZXsl::before{-webkit-transform:scale(var(--mdc-ripple-fg-scale,1));transform:scale(var(--mdc-ripple-fg-scale,1))}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d .VfPpkd-rymPhb-pZXsl::after{top:0;left:0;-webkit-transform:scale(0);transform:scale(0);-webkit-transform-origin:center center;transform-origin:center center}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-ZNMTqd .VfPpkd-rymPhb-pZXsl::after{top:var(--mdc-ripple-top,0);left:var(--mdc-ripple-left,0)}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-lJfZMc .VfPpkd-rymPhb-pZXsl::after{-webkit-animation:mdc-ripple-fg-radius-in 225ms forwards,mdc-ripple-fg-opacity-in 75ms forwards;animation:mdc-ripple-fg-radius-in 225ms forwards,mdc-ripple-fg-opacity-in 75ms forwards}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-Tv8l5d-OmS1vf .VfPpkd-rymPhb-pZXsl::after{-webkit-animation:mdc-ripple-fg-opacity-out .15s;animation:mdc-ripple-fg-opacity-out .15s;-webkit-transform:translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1));transform:translate(var(--mdc-ripple-fg-translate-end,0)) scale(var(--mdc-ripple-fg-scale,1))}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::before,:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::after{top:-50%;left:-50%;width:200%;height:200%}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d .VfPpkd-rymPhb-pZXsl::after{width:var(--mdc-ripple-fg-size,100%);height:var(--mdc-ripple-fg-size,100%)}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::before,:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::after{background-color:#000;background-color:var(--mdc-ripple-color,#000)}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b:hover .VfPpkd-rymPhb-pZXsl::before,:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-rymPhb-pZXsl::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-rymPhb-pZXsl::before,:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-rymPhb-pZXsl::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-rymPhb-pZXsl::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-rymPhb-pZXsl::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-press-opacity,.12)}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.12)}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-rymPhb-pZXsl::before{opacity:.12;opacity:var(--mdc-ripple-activated-opacity,.12)}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-rymPhb-pZXsl::before,:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-rymPhb-pZXsl::after{background-color:#6200ee;background-color:var(--mdc-ripple-color,var(--mdc-theme-primary,#6200ee))}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b:hover .VfPpkd-rymPhb-pZXsl::before,:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-rymPhb-pZXsl::before{opacity:.16;opacity:var(--mdc-ripple-hover-opacity,.16)}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-rymPhb-pZXsl::before,:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-rymPhb-pZXsl::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.24;opacity:var(--mdc-ripple-focus-opacity,.24)}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-rymPhb-pZXsl::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-rymPhb-pZXsl::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.24;opacity:var(--mdc-ripple-press-opacity,.24)}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.24)}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::before{opacity:.08;opacity:var(--mdc-ripple-selected-opacity,.08)}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::before,:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::after{background-color:#6200ee;background-color:var(--mdc-ripple-color,var(--mdc-theme-primary,#6200ee))}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-rymPhb-pZXsl::before,:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-rymPhb-pZXsl::before{opacity:.12;opacity:var(--mdc-ripple-hover-opacity,.12)}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-rymPhb-pZXsl::before,:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-rymPhb-pZXsl::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.2;opacity:var(--mdc-ripple-focus-opacity,.2)}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-rymPhb-pZXsl::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-rymPhb-pZXsl::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.2;opacity:var(--mdc-ripple-press-opacity,.2)}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.2)}:not(.VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me).VfPpkd-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl{position:relative;outline:none;overflow:hidden;position:absolute;top:0;left:0;width:100%;height:100%;pointer-events:none}.P2Hi5d,.mkMxfe,.OBi8lb,.P9QRxe,.vqjb4e,.y8Rdrf,.DMZ54e{font-family:Roboto,Arial,sans-serif;line-height:1.5rem;font-size:1rem;letter-spacing:.00625em;font-weight:400;color:#000;color:var(--mdc-theme-on-surface,#000)}.P2Hi5d .VfPpkd-StrnGf-rymPhb-IhFlZd,.mkMxfe .VfPpkd-StrnGf-rymPhb-IhFlZd,.OBi8lb .VfPpkd-StrnGf-rymPhb-IhFlZd,.P9QRxe .VfPpkd-StrnGf-rymPhb-IhFlZd,.vqjb4e .VfPpkd-StrnGf-rymPhb-IhFlZd,.y8Rdrf .VfPpkd-StrnGf-rymPhb-IhFlZd,.DMZ54e .VfPpkd-StrnGf-rymPhb-IhFlZd{color:rgb(95,99,104)}.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS{color:rgb(60,64,67)}.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c{opacity:.38}.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd,.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b{color:#000;color:var(--mdc-theme-on-surface,#000)}.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-f7MjDc,.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-f7MjDc,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-f7MjDc,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-f7MjDc,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-f7MjDc,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-f7MjDc,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-f7MjDc,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-f7MjDc,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-f7MjDc,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-f7MjDc,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-f7MjDc,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-f7MjDc,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-f7MjDc,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-f7MjDc{color:#000;color:var(--mdc-theme-on-surface,#000)}.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:0}.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd{background-color:rgb(232,240,254)}.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before,.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::after,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::after,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::after,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::after,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::after,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::after,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::after{background-color:rgb(26,115,232);background-color:var(--mdc-ripple-color,rgb(26,115,232))}.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before,.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before,.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}@media (-ms-high-contrast:active),screen and (forced-colors:active){.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS{color:GrayText}.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.OBi8lb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.P9QRxe .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.vqjb4e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.y8Rdrf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.DMZ54e .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c{opacity:1}}.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b{padding-left:24px;padding-right:16px}[dir=rtl] .P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b,.P2Hi5d .VfPpkd-StrnGf-rymPhb-ibnC6b[dir=rtl]{padding-left:16px;padding-right:24px}.P2Hi5d .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc{margin-left:24px;margin-right:0;width:calc(100% - 24px)}[dir=rtl] .P2Hi5d .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc,.P2Hi5d .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc[dir=rtl]{margin-left:0;margin-right:24px}.P2Hi5d .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg{width:calc(100% - 16px)}.P2Hi5d .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg{margin-left:24px;margin-right:0;width:calc(100% - 40px)}[dir=rtl] .P2Hi5d .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg,.P2Hi5d .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg[dir=rtl]{margin-left:0;margin-right:24px}.P2Hi5d .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2{margin-left:24px;margin-right:0;width:calc(100% - 24px)}[dir=rtl] .P2Hi5d .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2,.P2Hi5d .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2[dir=rtl]{margin-left:0;margin-right:24px}.P2Hi5d .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2{margin-left:24px;margin-right:0;width:calc(100% - 40px)}[dir=rtl] .P2Hi5d .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2,.P2Hi5d .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2[dir=rtl]{margin-left:0;margin-right:24px}.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-f7MjDc{margin-left:0;margin-right:16px}[dir=rtl] .mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-f7MjDc,.mkMxfe .VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-f7MjDc[dir=rtl]{margin-left:16px;margin-right:0}.mkMxfe .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc{margin-left:56px;margin-right:0;width:calc(100% - 56px)}[dir=rtl] .mkMxfe .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc,.mkMxfe .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc[dir=rtl]{margin-left:0;margin-right:56px}.mkMxfe .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg{width:calc(100% - 16px)}.mkMxfe .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg{margin-left:56px;margin-right:0;width:calc(100% - 72px)}[dir=rtl] .mkMxfe .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg,.mkMxfe .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg[dir=rtl]{margin-left:0;margin-right:56px}.mkMxfe .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2{margin-left:16px;margin-right:0;width:calc(100% - 16px)}[dir=rtl] .mkMxfe .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2,.mkMxfe .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-QFlW2[dir=rtl]{margin-left:0;margin-right:16px}.mkMxfe .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2{margin-left:16px;margin-right:0;width:calc(100% - 32px)}[dir=rtl] .mkMxfe .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2,.mkMxfe .VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-M1Soyc.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-UbuQg.VfPpkd-StrnGf-rymPhb-clz4Ic-OWXEXe-YbohUe-QFlW2[dir=rtl]{margin-left:0;margin-right:16px}.r6B9Fd{font-family:Roboto,Arial,sans-serif;line-height:1.5rem;font-size:1rem;letter-spacing:.00625em;font-weight:400}.r6B9Fd .VfPpkd-rymPhb-Gtdoyb,.r6B9Fd .VfPpkd-rymPhb-fpDzbe-fmcmS{color:rgb(60,64,67)}.r6B9Fd .VfPpkd-rymPhb-L8ivfd-fmcmS,.r6B9Fd .VfPpkd-rymPhb-bC5pod-fmcmS,.r6B9Fd .VfPpkd-rymPhb-JMEf7e{color:rgb(95,99,104)}.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb,.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e,.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-Gtdoyb,.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-fpDzbe-fmcmS,.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-L8ivfd-fmcmS,.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-bC5pod-fmcmS,.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb,.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e,.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e{color:rgb(60,64,67)}.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-KkROqb,.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-Gtdoyb,.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-JMEf7e{opacity:.38}.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-Gtdoyb,.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-fpDzbe-fmcmS,.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-rymPhb-Gtdoyb,.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-rymPhb-fpDzbe-fmcmS,.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb,.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb{color:rgb(60,64,67)}.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::before{opacity:0}.r6B9Fd .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd{background-color:rgb(232,240,254)}.r6B9Fd .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::before,.r6B9Fd .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::after{background-color:rgb(26,115,232);background-color:var(--mdc-ripple-color,rgb(26,115,232))}.r6B9Fd .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-rymPhb-pZXsl::before,.r6B9Fd .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-rymPhb-pZXsl::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.r6B9Fd .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-rymPhb-pZXsl::before,.r6B9Fd .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-rymPhb-pZXsl::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.r6B9Fd .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-rymPhb-pZXsl::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.r6B9Fd .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-rymPhb-pZXsl::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.r6B9Fd .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}@media screen and (forced-colors:active){.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-Gtdoyb,.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-fpDzbe-fmcmS,.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-L8ivfd-fmcmS,.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-bC5pod-fmcmS,.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb,.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e,.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e{color:GrayText}.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-KkROqb,.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-Gtdoyb,.r6B9Fd .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-JMEf7e{opacity:1}}.uTZ9Lb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-KkROqb,.FvXOfd.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-KkROqb,.QrsYgb.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-KkROqb,.gfwIBd.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-KkROqb{-webkit-align-self:center;align-self:center;margin-top:0}.HiC7Nc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc{height:56px}.HiC7Nc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-HiaYvf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc,.HiC7Nc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-aTv5jf.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-Woal0c-RWgCYc{height:72px}.UbEQCe.VfPpkd-rymPhb-ibnC6b{padding-left:0;padding-right:auto}[dir=rtl] .UbEQCe.VfPpkd-rymPhb-ibnC6b,.UbEQCe.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:auto;padding-right:0}.UbEQCe .VfPpkd-rymPhb-KkROqb{margin-left:16px;margin-right:16px}[dir=rtl] .UbEQCe .VfPpkd-rymPhb-KkROqb,.UbEQCe .VfPpkd-rymPhb-KkROqb[dir=rtl]{margin-left:16px;margin-right:16px}.rKASPc.VfPpkd-rymPhb-ibnC6b{padding-left:0;padding-right:auto}[dir=rtl] .rKASPc.VfPpkd-rymPhb-ibnC6b,.rKASPc.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:auto;padding-right:0}.rKASPc .VfPpkd-rymPhb-KkROqb{margin-left:8px;margin-right:8px}[dir=rtl] .rKASPc .VfPpkd-rymPhb-KkROqb,.rKASPc .VfPpkd-rymPhb-KkROqb[dir=rtl]{margin-left:8px;margin-right:8px}.rKASPc.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-KkROqb{-webkit-align-self:flex-start;align-self:flex-start;margin-top:8px}.U5k4Fd.VfPpkd-rymPhb-ibnC6b{padding-left:0;padding-right:auto}[dir=rtl] .U5k4Fd.VfPpkd-rymPhb-ibnC6b,.U5k4Fd.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:auto;padding-right:0}.U5k4Fd .VfPpkd-rymPhb-KkROqb{margin-left:8px;margin-right:8px}[dir=rtl] .U5k4Fd .VfPpkd-rymPhb-KkROqb,.U5k4Fd .VfPpkd-rymPhb-KkROqb[dir=rtl]{margin-left:8px;margin-right:8px}.U5k4Fd.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-KkROqb{-webkit-align-self:flex-start;align-self:flex-start;margin-top:8px}.ifEyr.VfPpkd-rymPhb-ibnC6b{padding-left:0;padding-right:auto}[dir=rtl] .ifEyr.VfPpkd-rymPhb-ibnC6b,.ifEyr.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:auto;padding-right:0}.ifEyr .VfPpkd-rymPhb-KkROqb{margin-left:8px;margin-right:8px}[dir=rtl] .ifEyr .VfPpkd-rymPhb-KkROqb,.ifEyr .VfPpkd-rymPhb-KkROqb[dir=rtl]{margin-left:8px;margin-right:8px}.ifEyr.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-aSi1db-MCEKJb .VfPpkd-rymPhb-KkROqb{-webkit-align-self:flex-start;align-self:flex-start;margin-top:8px}.SNowt.VfPpkd-rymPhb-ibnC6b{padding-left:auto;padding-right:0}[dir=rtl] .SNowt.VfPpkd-rymPhb-ibnC6b,.SNowt.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:0;padding-right:auto}.SNowt .VfPpkd-rymPhb-JMEf7e{margin-left:8px;margin-right:16px}[dir=rtl] .SNowt .VfPpkd-rymPhb-JMEf7e,.SNowt .VfPpkd-rymPhb-JMEf7e[dir=rtl]{margin-left:16px;margin-right:8px}.tfmWAf.VfPpkd-rymPhb-ibnC6b{padding-left:auto;padding-right:0}[dir=rtl] .tfmWAf.VfPpkd-rymPhb-ibnC6b,.tfmWAf.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:0;padding-right:auto}.tfmWAf .VfPpkd-rymPhb-JMEf7e{margin-left:8px;margin-right:16px}[dir=rtl] .tfmWAf .VfPpkd-rymPhb-JMEf7e,.tfmWAf .VfPpkd-rymPhb-JMEf7e[dir=rtl]{margin-left:16px;margin-right:8px}.axtYbd.VfPpkd-rymPhb-ibnC6b{padding-left:auto;padding-right:0}[dir=rtl] .axtYbd.VfPpkd-rymPhb-ibnC6b,.axtYbd.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:0;padding-right:auto}.axtYbd .VfPpkd-rymPhb-JMEf7e{margin-left:16px;margin-right:24px}[dir=rtl] .axtYbd .VfPpkd-rymPhb-JMEf7e,.axtYbd .VfPpkd-rymPhb-JMEf7e[dir=rtl]{margin-left:24px;margin-right:16px}.aopLEb.VfPpkd-rymPhb-ibnC6b{padding-left:auto;padding-right:0}[dir=rtl] .aopLEb.VfPpkd-rymPhb-ibnC6b,.aopLEb.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:0;padding-right:auto}.aopLEb .VfPpkd-rymPhb-JMEf7e{margin-left:16px;margin-right:24px}[dir=rtl] .aopLEb .VfPpkd-rymPhb-JMEf7e,.aopLEb .VfPpkd-rymPhb-JMEf7e[dir=rtl]{margin-left:24px;margin-right:16px}.zlqiud.VfPpkd-rymPhb-ibnC6b{padding-left:auto;padding-right:0}[dir=rtl] .zlqiud.VfPpkd-rymPhb-ibnC6b,.zlqiud.VfPpkd-rymPhb-ibnC6b[dir=rtl]{padding-left:0;padding-right:auto}.zlqiud .VfPpkd-rymPhb-JMEf7e{margin-left:16px;margin-right:24px}[dir=rtl] .zlqiud .VfPpkd-rymPhb-JMEf7e,.zlqiud .VfPpkd-rymPhb-JMEf7e[dir=rtl]{margin-left:24px;margin-right:16px}.isC8Y.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe{padding-left:24px;padding-right:auto}[dir=rtl] .isC8Y.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe,.isC8Y.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-M1Soyc-YbohUe[dir=rtl]{padding-left:auto;padding-right:24px}.MCs1Pd{padding-left:24px;padding-right:24px}[dir=rtl] .MCs1Pd,.MCs1Pd[dir=rtl]{padding-left:24px;padding-right:24px}.e6pQl.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe{padding-left:auto;padding-right:24px}[dir=rtl] .e6pQl.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe,.e6pQl.VfPpkd-rymPhb-clz4Ic-OWXEXe-SfQLQb-UbuQg-YbohUe[dir=rtl]{padding-left:24px;padding-right:auto}[dir=rtl] .e6pQl,.e6pQl[dir=rtl]{padding:0}.VfPpkd-xl07Ob-XxIAqe{display:none;position:absolute;box-sizing:border-box;margin:0;padding:0;-webkit-transform:scale(1);transform:scale(1);-webkit-transform-origin:top left;transform-origin:top left;opacity:0;overflow:auto;will-change:transform,opacity;box-shadow:0 5px 5px -3px rgba(0,0,0,.2),0 8px 10px 1px rgba(0,0,0,.14),0 3px 14px 2px rgba(0,0,0,.12);transform-origin-left:top left;transform-origin-right:top right}.VfPpkd-xl07Ob-XxIAqe:focus{outline:none}.VfPpkd-xl07Ob-XxIAqe-OWXEXe-oT9UPb-FNFY6c{display:inline-block;-webkit-transform:scale(.8);transform:scale(.8);opacity:0}.VfPpkd-xl07Ob-XxIAqe-OWXEXe-FNFY6c{display:inline-block;-webkit-transform:scale(1);transform:scale(1);opacity:1}.VfPpkd-xl07Ob-XxIAqe-OWXEXe-oT9UPb-xTMeO{display:inline-block;opacity:0}[dir=rtl] .VfPpkd-xl07Ob-XxIAqe,.VfPpkd-xl07Ob-XxIAqe[dir=rtl]{transform-origin-left:top right;transform-origin-right:top left}.VfPpkd-xl07Ob-XxIAqe-OWXEXe-oYxtQd{position:relative;overflow:visible}.VfPpkd-xl07Ob-XxIAqe-OWXEXe-qbOKL{position:fixed}.VfPpkd-xl07Ob-XxIAqe-OWXEXe-tsQazb{width:100%}.VfPpkd-xl07Ob-XxIAqe{max-width:calc(100vw - 32px);max-width:var(--mdc-menu-max-width,calc(100vw - 32px));max-height:calc(100vh - 32px);max-height:var(--mdc-menu-max-height,calc(100vh - 32px));z-index:8;-webkit-transition:opacity .03s linear,height .25s cubic-bezier(0,0,.2,1),-webkit-transform .12s cubic-bezier(0,0,.2,1);transition:opacity .03s linear,height .25s cubic-bezier(0,0,.2,1),-webkit-transform .12s cubic-bezier(0,0,.2,1);transition:opacity .03s linear,transform .12s cubic-bezier(0,0,.2,1),height .25s cubic-bezier(0,0,.2,1);transition:opacity .03s linear,transform .12s cubic-bezier(0,0,.2,1),height .25s cubic-bezier(0,0,.2,1),-webkit-transform .12s cubic-bezier(0,0,.2,1);background-color:#fff;background-color:var(--mdc-theme-surface,#fff);color:#000;color:var(--mdc-theme-on-surface,#000);border-radius:4px;border-radius:var(--mdc-shape-medium,4px)}.VfPpkd-xl07Ob-XxIAqe-OWXEXe-oT9UPb-xTMeO{-webkit-transition:opacity 75ms linear;transition:opacity 75ms linear}.UQ5E0{box-shadow:0 3px 5px -1px rgba(0,0,0,.2),0 6px 10px 0 rgba(0,0,0,.14),0 1px 18px 0 rgba(0,0,0,.12)}.VfPpkd-xl07Ob{min-width:112px;min-width:var(--mdc-menu-min-width,112px)}.VfPpkd-xl07Ob .VfPpkd-StrnGf-rymPhb-IhFlZd,.VfPpkd-xl07Ob .VfPpkd-StrnGf-rymPhb-f7MjDc{color:rgba(0,0,0,.87)}.VfPpkd-xl07Ob .VfPpkd-xl07Ob-ibnC6b-OWXEXe-eKm5Fc-FNFY6c .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:.04}.VfPpkd-xl07Ob .VfPpkd-xl07Ob-ibnC6b-OWXEXe-eKm5Fc-FNFY6c .VfPpkd-rymPhb-pZXsl::before{opacity:.04}.VfPpkd-xl07Ob .VfPpkd-StrnGf-rymPhb{color:rgba(0,0,0,.87)}.VfPpkd-xl07Ob .VfPpkd-StrnGf-rymPhb,.VfPpkd-xl07Ob .VfPpkd-rymPhb{position:relative;border-radius:inherit}.VfPpkd-xl07Ob .VfPpkd-StrnGf-rymPhb .VfPpkd-BFbNVe-bF1uUb,.VfPpkd-xl07Ob .VfPpkd-rymPhb .VfPpkd-BFbNVe-bF1uUb{width:100%;height:100%;top:0;left:0}.VfPpkd-xl07Ob .VfPpkd-StrnGf-rymPhb::before,.VfPpkd-xl07Ob .VfPpkd-rymPhb::before{position:absolute;box-sizing:border-box;width:100%;height:100%;top:0;left:0;border:1px solid transparent;border-radius:inherit;content:"";pointer-events:none}@media screen and (forced-colors:active){.VfPpkd-xl07Ob .VfPpkd-StrnGf-rymPhb::before,.VfPpkd-xl07Ob .VfPpkd-rymPhb::before{border-color:CanvasText}}.VfPpkd-xl07Ob .VfPpkd-StrnGf-rymPhb-clz4Ic{margin:8px 0}.VfPpkd-xl07Ob .VfPpkd-StrnGf-rymPhb-ibnC6b{-webkit-user-select:none;user-select:none}.VfPpkd-xl07Ob .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me{cursor:auto}.VfPpkd-xl07Ob a.VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-b9t22c,.VfPpkd-xl07Ob a.VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-f7MjDc{pointer-events:none}.VfPpkd-qPzbhe-JNdkSc{padding:0;fill:currentColor}.VfPpkd-qPzbhe-JNdkSc .VfPpkd-StrnGf-rymPhb-ibnC6b{padding-left:56px;padding-right:16px}[dir=rtl] .VfPpkd-qPzbhe-JNdkSc .VfPpkd-StrnGf-rymPhb-ibnC6b,.VfPpkd-qPzbhe-JNdkSc .VfPpkd-StrnGf-rymPhb-ibnC6b[dir=rtl]{padding-left:16px;padding-right:56px}.VfPpkd-qPzbhe-JNdkSc .VfPpkd-qPzbhe-JNdkSc-Bz112c{left:16px;right:auto;visibility:hidden;position:absolute;top:50%;-webkit-transform:translateY(-50%);transform:translateY(-50%);-webkit-transition-property:visibility;transition-property:visibility;-webkit-transition-delay:75ms;transition-delay:75ms}[dir=rtl] .VfPpkd-qPzbhe-JNdkSc .VfPpkd-qPzbhe-JNdkSc-Bz112c,.VfPpkd-qPzbhe-JNdkSc .VfPpkd-qPzbhe-JNdkSc-Bz112c[dir=rtl]{left:auto;right:16px}.VfPpkd-xl07Ob-ibnC6b-OWXEXe-gk6SMd .VfPpkd-qPzbhe-JNdkSc-Bz112c{display:inline;visibility:visible}.q6oraf{box-shadow:0 3px 5px -1px rgba(0,0,0,.2),0 6px 10px 0 rgba(0,0,0,.14),0 1px 18px 0 rgba(0,0,0,.12)}.q6oraf .VfPpkd-StrnGf-rymPhb{font-family:Roboto,Arial,sans-serif;line-height:1.5rem;font-size:1rem;letter-spacing:.00625em;font-weight:400;color:#000;color:var(--mdc-theme-on-surface,#000)}.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-IhFlZd{color:rgb(95,99,104)}.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS{color:rgb(60,64,67)}.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c{opacity:.38}.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd,.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b{color:#000;color:var(--mdc-theme-on-surface,#000)}.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-f7MjDc,.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-f7MjDc{color:#000;color:var(--mdc-theme-on-surface,#000)}.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:0}.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd{background-color:rgb(232,240,254)}.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before,.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::after{background-color:rgb(26,115,232);background-color:var(--mdc-ripple-color,rgb(26,115,232))}.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before,.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before,.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}@media (-ms-high-contrast:active),screen and (forced-colors:active){.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS{color:GrayText}.q6oraf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c{opacity:1}}.FliLIb{box-sizing:border-box;display:inline-block}.FliLIb .u3bW4e{box-shadow:0px 6px 10px 0px rgba(0,0,0,.14),0px 1px 18px 0px rgba(0,0,0,.12),0px 3px 5px -1px rgba(0,0,0,.2)}.FliLIb.eLNT1d{display:none}.FliLIb .q6oraf .VfPpkd-rymPhb,.FliLIb .ksBjEc{font-size:inherit}.FliLIb .TrZEUc .WpHeLc{position:absolute}.FliLIb .qIypjc:not(:disabled){color:#fff}.xYnMae .VfPpkd-Jh9lGc{box-sizing:content-box}.uRo0Xe .snByac{font-weight:500;line-height:1.4286}.FliLIb .uRo0Xe{min-width:0}.uRo0Xe .snByac{margin:8px 8px;text-transform:none}.stUf5b.WS4XDd{border:0;max-height:1.3333333em;padding:0 2px;vertical-align:middle;width:auto}.G5XIyb{border:0;object-fit:contain}.G5XIyb.WS4XDd{border:0;max-height:1.3333333em;padding:0 2px;vertical-align:middle;width:auto}.YZrg6{-webkit-box-align:center;-webkit-align-items:center;align-items:center;background:#fff;border:1px solid rgb(218,220,224);box-sizing:border-box;color:rgb(60,64,67);cursor:pointer;display:-webkit-inline-box;display:-webkit-inline-flex;display:inline-flex;font-family:"Google Sans","Noto Sans Myanmar UI",arial,sans-serif;font-size:14px;font-weight:500;letter-spacing:.25px;max-width:100%;position:relative}.YZrg6::after{bottom:-1px;border:1px solid transparent;content:"";left:-1px;position:absolute;right:-1px;top:-1px}.YZrg6:focus,.YZrg6.u3bW4e{background:rgba(60,64,67,0.122);outline:none}.YZrg6:focus-visible::after{bottom:-5px;border:2px solid rgb(24,90,188);border-radius:20px;box-shadow:0 0 0 2px rgb(232,240,254);content:"";left:-5px;position:absolute;right:-5px;top:-5px}.YZrg6:hover:not(:focus-visible)::after{background:rgba(60,64,67,0.039)}.YZrg6:focus:not(:focus-visible)::after,.YZrg6:hover:not(:focus-visible)::after,.YZrg6.u3bW4e{border-color:rgb(218,220,224)}.YZrg6.qs41qe{color:rgb(60,64,67)}.YZrg6.qs41qe:not(:focus-visible)::after{background:rgba(60,64,67,0.122);border-color:rgb(60,64,67)}.SOOv2c{color:rgb(26,115,232);font-size:12px}.HnRr5d{border-radius:16px;padding:0 15px 0 15px}.HnRr5d.SOOv2c{border-radius:12px;padding:0 10px 0 10px}.HnRr5d.iiFyne{padding-right:7px}.HnRr5d.cd29Sd{padding-left:5px}.HnRr5d.SOOv2c.iiFyne{padding-right:7px}.HnRr5d.SOOv2c.cd29Sd{padding-left:2px}.HnRr5d::after{border-radius:16px}.HnRr5d.SOOv2c::after{border-radius:12px}.gPHLDe{border-radius:10px;height:20px;margin-right:8px}.gPHLDe .stUf5b,.gPHLDe .G5XIyb{border-radius:50%;color:rgb(60,64,67);display:block;height:20px;width:20px}.KTeGk{direction:ltr;text-align:left;overflow:hidden;text-overflow:ellipsis;white-space:nowrap}.HnRr5d .KTeGk{line-height:30px}.HnRr5d.SOOv2c .KTeGk{line-height:22px}.krLnGe{color:rgb(60,64,67);-webkit-flex-shrink:0;flex-shrink:0;height:18px;margin-left:4px;-webkit-transition:-webkit-transform .2s cubic-bezier(.4,0,.2,1);transition:-webkit-transform .2s cubic-bezier(.4,0,.2,1);transition:transform .2s cubic-bezier(.4,0,.2,1);transition:transform .2s cubic-bezier(.4,0,.2,1),-webkit-transform .2s cubic-bezier(.4,0,.2,1);width:18px}.YZrg6.sMVRZe .krLnGe{-webkit-transform:rotate(180deg);transform:rotate(180deg)}.SOOv2c .krLnGe{height:16px;width:16px}.MSBt4d{display:block;height:100%;width:100%}.aTzEhb{margin:16px 0;outline:none}.aTzEhb+.aTzEhb{margin-top:24px}.aTzEhb:first-child{margin-top:0}.aTzEhb:last-child{margin-bottom:0}.AORPd{-webkit-border-radius:8px;border-radius:8px;padding:16px}.AORPd>:first-child{margin-top:0}.AORPd>:last-child{margin-bottom:0}.AORPd .kV95Wc{color:rgb(32,33,36)}.AORPd .CxRgyd{color:rgb(32,33,36)}.AORPd.YFdWic .CxRgyd{color:rgb(95,99,104);margin-top:4px;padding:0}.AORPd.YFdWic .IdEPtc,.AORPd.YFdWic .CxRgyd{margin-left:64px;width:-webkit-calc(100% - 64px);width:calc(100% - 64px)}.AORPd.YFdWic:not(.S7S4N) .IdEPtc{margin-left:0;width:0}.AORPd:not(.S7S4N)>.CxRgyd{margin-top:0}.AORPd.sj692e{background:rgb(232,240,254)}.AORPd.Xq8bDe{background:rgb(252,232,230)}.AORPd.rNe0id{background:rgb(254,247,224)}.AORPd.YFdWic{border:1px solid rgb(218,220,224);-webkit-box-sizing:border-box;box-sizing:border-box;min-height:80px;position:relative}.AORPd:not(.S7S4N){display:-webkit-box;display:-webkit-flex;display:-webkit-box;display:-webkit-flex;display:flex}.aTzEhb.eLNT1d{display:none}.aTzEhb.RDPZE{opacity:.5;pointer-events:none}.aTzEhb.RDPZE .aTzEhb.RDPZE{opacity:1}.wfep7d{border:1px solid rgb(218,220,224);-webkit-border-radius:8px;border-radius:8px;padding:16px}.wfep7d .UST9Bf{display:-webkit-box;display:-webkit-flex;display:-webkit-box;display:-webkit-flex;display:flex;-webkit-box-pack:end;-webkit-justify-content:flex-end;-webkit-justify-content:flex-end;justify-content:flex-end;margin-top:16px}.wfep7d .UST9Bf .xYnMae{margin-bottom:0;margin-top:0}.vEFDtd{border-bottom:1px solid rgb(218,220,224);display:-webkit-box;display:-webkit-flex;display:-webkit-box;display:-webkit-flex;display:flex;-webkit-box-orient:vertical;-webkit-box-direction:normal;-webkit-flex-direction:column;-webkit-flex-direction:column;flex-direction:column}.vEFDtd .V9RXW .rBUW7e,.vEFDtd .vEFDtd:last-child{border-bottom:0}.vEFDtd .vEFDtd:last-child .L9iFZc{padding-bottom:0}.vEFDtd.D6kf4b{border-bottom:0}.IdEPtc:empty,.yMb59d:empty{display:none}.IdEPtc>:first-child{margin-top:0;padding-top:0}.IdEPtc>:last-child{margin-bottom:0;padding-bottom:0}.UWVyoc{margin:0 0 8px}.vEFDtd[data-expand-type="1"] .L9iFZc,.aTzEhb[data-expand-type="1"] .A6OHve{cursor:pointer}.vEFDtd .L9iFZc{padding-bottom:16px}.kV95Wc{-webkit-box-align:center;-webkit-align-items:center;-webkit-align-items:center;align-items:center;color:rgb(32,33,36);display:-webkit-box;display:-webkit-flex;display:-webkit-box;display:-webkit-flex;display:flex;font-family:"Google Sans","Noto Sans Myanmar UI",arial,sans-serif;font-size:16px;font-weight:500;letter-spacing:.1px;line-height:1.5;margin-top:0;margin-bottom:0;padding:0}.vEFDtd.u3bW4e .kV95Wc{position:relative}.vEFDtd[data-expand-type="1"].u3bW4e .kV95Wc::after{background:rgba(26,115,232,0.149);-webkit-border-radius:8px;border-radius:8px;bottom:-4px;content:"";left:-8px;position:absolute;right:-8px;top:-4px;z-index:-1}.A6OHve{background:none;border:none;color:inherit;-webkit-box-flex:1;-webkit-flex-grow:1;-webkit-box-flex:1;box-flex:1;-webkit-flex-grow:1;flex-grow:1;font:inherit;margin:0;outline:0;padding:0;text-align:inherit}.A6OHve::-moz-focus-inner{border:0}.A6OHve [jsslot]{position:relative}.jhXB3b{margin-left:16px}.jhXB3b .Z6O26d{-webkit-box-align:center;-webkit-align-items:center;-webkit-align-items:center;align-items:center;display:-webkit-box;display:-webkit-flex;display:-webkit-box;display:-webkit-flex;display:flex;height:24px;-webkit-box-pack:center;-webkit-justify-content:center;-webkit-justify-content:center;justify-content:center;-webkit-transition:-webkit-transform .2s cubic-bezier(0.4,0,0.2,1);-webkit-transition:-webkit-transform .2s cubic-bezier(0.4,0,0.2,1);transition:-webkit-transform .2s cubic-bezier(0.4,0,0.2,1);-webkit-transition:transform .2s cubic-bezier(0.4,0,0.2,1);transition:transform .2s cubic-bezier(0.4,0,0.2,1);-webkit-transition:transform .2s cubic-bezier(0.4,0,0.2,1),-webkit-transform .2s cubic-bezier(0.4,0,0.2,1);transition:transform .2s cubic-bezier(0.4,0,0.2,1),-webkit-transform .2s cubic-bezier(0.4,0,0.2,1);width:24px}.vEFDtd .jhXB3b,.vEFDtd .A6OHve,.vEFDtd .yiP64c{pointer-events:none}.vEFDtd.jVwmLb .Z6O26d{-webkit-transform:rotate(-180deg);-webkit-transform:rotate(-180deg);transform:rotate(-180deg)}.yiP64c{color:rgb(95,99,104);-webkit-flex-shrink:0;-webkit-flex-shrink:0;flex-shrink:0;height:20px;margin-right:16px;width:20px}.yiP64c .d7Plee{height:100%;width:100%}.AORPd .yiP64c{margin-top:0}.AORPd.sj692e .yiP64c{color:rgb(25,103,210)}.AORPd.Xq8bDe .yiP64c{color:rgb(197,34,31)}.AORPd.rNe0id .yiP64c{color:rgb(234,134,0)}.AORPd.YFdWic .yiP64c{height:48px;left:16px;position:absolute;top:16px;width:48px}.yMb59d{color:rgb(95,99,104);font-size:14px;font-weight:400;line-height:1.4286;margin-top:8px}.CxRgyd{margin:auto -24px;padding-left:24px;padding-right:24px;margin-bottom:16px;margin-top:10px}@media (min-width:450px){.CxRgyd{margin:auto -40px;padding-left:40px;padding-right:40px;margin-bottom:16px;margin-top:10px}}.wfep7d .CxRgyd{margin-bottom:0;margin-top:16px}.IdEPtc:empty+.CxRgyd{margin-top:0}.CxRgyd:only-child{margin-bottom:0;margin-top:0}.vEFDtd .CxRgyd{margin-top:0;overflow-y:hidden;-webkit-transition:.2s cubic-bezier(0.4,0,0.2,1);-webkit-transition:.2s cubic-bezier(0.4,0,0.2,1);transition:.2s cubic-bezier(0.4,0,0.2,1)}.vEFDtd.jVwmLb .CxRgyd{margin-bottom:0;margin-top:0;max-height:0;opacity:0;visibility:hidden}.CxRgyd>[jsslot]>:first-child:not(section){margin-top:0;padding-top:0}.CxRgyd>[jsslot]>:last-child:not(section){margin-bottom:0;padding-bottom:0}.w7wqLd{-webkit-align-self:center;-webkit-align-self:center;align-self:center;margin-bottom:0}.x3iGMd{border-bottom:1px solid rgb(218,220,224);display:-webkit-box;display:-webkit-flex;display:-webkit-box;display:-webkit-flex;display:flex;-webkit-box-orient:horizontal;-webkit-box-direction:normal;-webkit-flex-direction:row;-webkit-flex-direction:row;flex-direction:row;-webkit-box-pack:center;-webkit-justify-content:center;-webkit-justify-content:center;justify-content:center;height:0;margin-bottom:24px;margin-top:12px}.aQPcpb{background:#fff;display:-webkit-box;display:-webkit-flex;display:-webkit-box;display:-webkit-flex;display:flex;height:24px;margin-top:-12px}.D6kf4b:not(.jVwmLb) .x3iGMd{display:none}.D6kf4b .VBGMK:focus-visible{outline:none;position:relative}.D6kf4b .VBGMK:focus-visible::after{border:2px solid #185abc;border-radius:6px;bottom:0;box-shadow:0 0 0 2px #e8f0fe;content:"";left:0;position:absolute;right:0;top:0}.VfPpkd-Sx9Kwc .VfPpkd-P5QLlc{background-color:#fff;background-color:var(--mdc-theme-surface,#fff)}.VfPpkd-Sx9Kwc .VfPpkd-IE5DDf,.VfPpkd-Sx9Kwc .VfPpkd-P5QLlc-GGAcbc{background-color:rgba(0,0,0,.32)}.VfPpkd-Sx9Kwc .VfPpkd-k2Wrsb{color:rgba(0,0,0,.87)}.VfPpkd-Sx9Kwc .VfPpkd-cnG4Wd{color:rgba(0,0,0,.6)}.VfPpkd-Sx9Kwc .VfPpkd-zMU9ub{color:#000;color:var(--mdc-theme-on-surface,#000)}.VfPpkd-Sx9Kwc .VfPpkd-zMU9ub .VfPpkd-Bz112c-Jh9lGc::before,.VfPpkd-Sx9Kwc .VfPpkd-zMU9ub .VfPpkd-Bz112c-Jh9lGc::after{background-color:#000;background-color:var(--mdc-ripple-color,var(--mdc-theme-on-surface,#000))}.VfPpkd-Sx9Kwc .VfPpkd-zMU9ub:hover .VfPpkd-Bz112c-Jh9lGc::before,.VfPpkd-Sx9Kwc .VfPpkd-zMU9ub.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Bz112c-Jh9lGc::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.VfPpkd-Sx9Kwc .VfPpkd-zMU9ub.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Bz112c-Jh9lGc::before,.VfPpkd-Sx9Kwc .VfPpkd-zMU9ub:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Bz112c-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.VfPpkd-Sx9Kwc .VfPpkd-zMU9ub:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Bz112c-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.VfPpkd-Sx9Kwc .VfPpkd-zMU9ub:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Bz112c-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-press-opacity,.12)}.VfPpkd-Sx9Kwc .VfPpkd-zMU9ub.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.12)}.VfPpkd-Sx9Kwc.VfPpkd-Sx9Kwc-OWXEXe-s2gQvd .VfPpkd-k2Wrsb,.VfPpkd-Sx9Kwc.VfPpkd-Sx9Kwc-OWXEXe-s2gQvd .VfPpkd-T0kwCb,.VfPpkd-Sx9Kwc.VfPpkd-Sx9Kwc-OWXEXe-s2gQvd.VfPpkd-Sx9Kwc-XuHpsb-clz4Ic-yePe5c .VfPpkd-T0kwCb{border-color:rgba(0,0,0,.12)}.VfPpkd-Sx9Kwc.VfPpkd-Sx9Kwc-OWXEXe-s2gQvd .VfPpkd-k2Wrsb{border-bottom:1px solid rgba(0,0,0,.12);margin-bottom:0}.VfPpkd-Sx9Kwc.VfPpkd-Sx9Kwc-XuHpsb-clz4Ic-tJHJj.VfPpkd-Sx9Kwc-OWXEXe-n9oEIb .VfPpkd-oclYLd{box-shadow:0 3px 1px -2px rgba(0,0,0,.2),0 2px 2px 0 rgba(0,0,0,.14),0 1px 5px 0 rgba(0,0,0,.12)}.VfPpkd-Sx9Kwc .VfPpkd-P5QLlc{border-radius:4px;border-radius:var(--mdc-shape-medium,4px)}.VfPpkd-P5QLlc{box-shadow:0 11px 15px -7px rgba(0,0,0,.2),0 24px 38px 3px rgba(0,0,0,.14),0 9px 46px 8px rgba(0,0,0,.12)}.VfPpkd-k2Wrsb{-moz-osx-font-smoothing:grayscale;-webkit-font-smoothing:antialiased;font-family:Roboto,sans-serif;font-family:var(--mdc-typography-headline6-font-family,var(--mdc-typography-font-family,Roboto,sans-serif));font-size:1.25rem;font-size:var(--mdc-typography-headline6-font-size,1.25rem);line-height:2rem;line-height:var(--mdc-typography-headline6-line-height,2rem);font-weight:500;font-weight:var(--mdc-typography-headline6-font-weight,500);letter-spacing:.0125em;letter-spacing:var(--mdc-typography-headline6-letter-spacing,.0125em);text-decoration:inherit;-webkit-text-decoration:var(--mdc-typography-headline6-text-decoration,inherit);text-decoration:var(--mdc-typography-headline6-text-decoration,inherit);text-transform:inherit;text-transform:var(--mdc-typography-headline6-text-transform,inherit)}.VfPpkd-cnG4Wd{-moz-osx-font-smoothing:grayscale;-webkit-font-smoothing:antialiased;font-family:Roboto,sans-serif;font-family:var(--mdc-typography-body1-font-family,var(--mdc-typography-font-family,Roboto,sans-serif));font-size:1rem;font-size:var(--mdc-typography-body1-font-size,1rem);line-height:1.5rem;line-height:var(--mdc-typography-body1-line-height,1.5rem);font-weight:400;font-weight:var(--mdc-typography-body1-font-weight,400);letter-spacing:.03125em;letter-spacing:var(--mdc-typography-body1-letter-spacing,.03125em);text-decoration:inherit;-webkit-text-decoration:var(--mdc-typography-body1-text-decoration,inherit);text-decoration:var(--mdc-typography-body1-text-decoration,inherit);text-transform:inherit;text-transform:var(--mdc-typography-body1-text-transform,inherit)}.VfPpkd-Sx9Kwc,.VfPpkd-IE5DDf{position:fixed;top:0;left:0;-webkit-box-align:center;-webkit-align-items:center;align-items:center;-webkit-box-pack:center;-webkit-justify-content:center;justify-content:center;box-sizing:border-box;width:100%;height:100%}.VfPpkd-Sx9Kwc{display:none;z-index:7;z-index:var(--mdc-dialog-z-index,7)}.VfPpkd-Sx9Kwc .VfPpkd-cnG4Wd{padding:20px 24px 20px 24px}.VfPpkd-Sx9Kwc .VfPpkd-P5QLlc{min-width:280px}@media (max-width:592px){.VfPpkd-Sx9Kwc .VfPpkd-P5QLlc{max-width:calc(100vw - 32px)}}@media (min-width:592px){.VfPpkd-Sx9Kwc .VfPpkd-P5QLlc{max-width:560px}}.VfPpkd-Sx9Kwc .VfPpkd-P5QLlc{max-height:calc(100% - 32px)}.VfPpkd-Sx9Kwc.VfPpkd-Sx9Kwc-OWXEXe-n9oEIb .VfPpkd-P5QLlc{max-width:none}@media (max-width:960px){.VfPpkd-Sx9Kwc.VfPpkd-Sx9Kwc-OWXEXe-n9oEIb .VfPpkd-P5QLlc{max-height:560px;width:560px}.VfPpkd-Sx9Kwc.VfPpkd-Sx9Kwc-OWXEXe-n9oEIb .VfPpkd-P5QLlc .VfPpkd-zMU9ub-suEOdc-sM5MNb{position:relative;right:-12px}}@media (max-width:720px) and (max-width:672px){.VfPpkd-Sx9Kwc.VfPpkd-Sx9Kwc-OWXEXe-n9oEIb .VfPpkd-P5QLlc{width:calc(100vw - 112px)}}@media (max-width:720px) and (min-width:672px){.VfPpkd-Sx9Kwc.VfPpkd-Sx9Kwc-OWXEXe-n9oEIb .VfPpkd-P5QLlc{width:560px}}@media (max-width:720px) and (max-height:720px){.VfPpkd-Sx9Kwc.VfPpkd-Sx9Kwc-OWXEXe-n9oEIb .VfPpkd-P5QLlc{max-height:calc(100vh - 160px)}}@media (max-width:720px) and (min-height:720px){.VfPpkd-Sx9Kwc.VfPpkd-Sx9Kwc-OWXEXe-n9oEIb .VfPpkd-P5QLlc{max-height:560px}}@media (max-width:720px){.VfPpkd-Sx9Kwc.VfPpkd-Sx9Kwc-OWXEXe-n9oEIb .VfPpkd-P5QLlc .VfPpkd-zMU9ub-suEOdc-sM5MNb{position:relative;right:-12px}}@media (max-width:600px),(max-width:720px) and (max-height:400px),(min-width:720px) and (max-height:400px){.VfPpkd-Sx9Kwc.VfPpkd-Sx9Kwc-OWXEXe-n9oEIb .VfPpkd-P5QLlc{height:100%;max-height:100vh;max-width:100vw;width:100vw;border-radius:0}.VfPpkd-Sx9Kwc.VfPpkd-Sx9Kwc-OWXEXe-n9oEIb .VfPpkd-P5QLlc .VfPpkd-zMU9ub-suEOdc-sM5MNb{position:relative;-webkit-box-ordinal-group:0;-webkit-order:-1;order:-1;left:-12px}.VfPpkd-Sx9Kwc.VfPpkd-Sx9Kwc-OWXEXe-n9oEIb .VfPpkd-P5QLlc .VfPpkd-oclYLd{padding:0 16px 9px;-webkit-box-pack:start;-webkit-justify-content:flex-start;justify-content:flex-start}.VfPpkd-Sx9Kwc.VfPpkd-Sx9Kwc-OWXEXe-n9oEIb .VfPpkd-P5QLlc .VfPpkd-k2Wrsb{margin-left:-8px}}@media (min-width:960px){.VfPpkd-Sx9Kwc.VfPpkd-Sx9Kwc-OWXEXe-n9oEIb .VfPpkd-P5QLlc{width:calc(100vw - 400px)}.VfPpkd-Sx9Kwc.VfPpkd-Sx9Kwc-OWXEXe-n9oEIb .VfPpkd-P5QLlc .VfPpkd-zMU9ub-suEOdc-sM5MNb{position:relative;right:-12px}}.VfPpkd-Sx9Kwc.VfPpkd-IE5DDf-OWXEXe-L6cTce .VfPpkd-IE5DDf{opacity:0}.VfPpkd-IE5DDf{opacity:0;z-index:-1}.VfPpkd-wzTsW{display:-webkit-box;display:-webkit-flex;display:flex;-webkit-box-orient:horizontal;-webkit-box-direction:normal;-webkit-flex-direction:row;flex-direction:row;-webkit-box-align:center;-webkit-align-items:center;align-items:center;-webkit-justify-content:space-around;justify-content:space-around;box-sizing:border-box;height:100%;opacity:0;pointer-events:none}.VfPpkd-P5QLlc{position:relative;display:-webkit-box;display:-webkit-flex;display:flex;-webkit-box-orient:vertical;-webkit-box-direction:normal;-webkit-flex-direction:column;flex-direction:column;-webkit-box-flex:0;-webkit-flex-grow:0;flex-grow:0;-webkit-flex-shrink:0;flex-shrink:0;box-sizing:border-box;max-width:100%;max-height:100%;pointer-events:auto;overflow-y:auto;outline:0;-webkit-transform:scale(.8);transform:scale(.8)}.VfPpkd-P5QLlc .VfPpkd-BFbNVe-bF1uUb{width:100%;height:100%;top:0;left:0}[dir=rtl] .VfPpkd-P5QLlc,.VfPpkd-P5QLlc[dir=rtl]{text-align:right}@media (-ms-high-contrast:active),screen and (forced-colors:active){.VfPpkd-P5QLlc{outline:2px solid windowText}}.VfPpkd-P5QLlc::before{position:absolute;box-sizing:border-box;width:100%;height:100%;top:0;left:0;border:2px solid transparent;border-radius:inherit;content:"";pointer-events:none}@media screen and (forced-colors:active){.VfPpkd-P5QLlc::before{border-color:CanvasText}}@media screen and (-ms-high-contrast:active),screen and (-ms-high-contrast:none){.VfPpkd-P5QLlc::before{content:none}}.VfPpkd-k2Wrsb{display:block;margin-top:0;position:relative;-webkit-flex-shrink:0;flex-shrink:0;box-sizing:border-box;margin:0 0 1px;padding:0 24px 9px}.VfPpkd-k2Wrsb::before{display:inline-block;width:0;height:40px;content:"";vertical-align:0}[dir=rtl] .VfPpkd-k2Wrsb,.VfPpkd-k2Wrsb[dir=rtl]{text-align:right}.VfPpkd-Sx9Kwc-OWXEXe-s2gQvd .VfPpkd-k2Wrsb{margin-bottom:1px;padding-bottom:15px}.VfPpkd-Sx9Kwc-OWXEXe-n9oEIb .VfPpkd-oclYLd{-webkit-box-align:baseline;-webkit-align-items:baseline;align-items:baseline;border-bottom:1px solid transparent;display:-webkit-inline-box;display:-webkit-inline-flex;display:inline-flex;-webkit-box-pack:justify;-webkit-justify-content:space-between;justify-content:space-between;padding:0 24px 9px;z-index:1}@media screen and (forced-colors:active){.VfPpkd-Sx9Kwc-OWXEXe-n9oEIb .VfPpkd-oclYLd{border-bottom-color:CanvasText}}.VfPpkd-Sx9Kwc-OWXEXe-n9oEIb .VfPpkd-oclYLd .VfPpkd-zMU9ub-suEOdc-sM5MNb{position:relative;right:-12px}.VfPpkd-Sx9Kwc-OWXEXe-n9oEIb .VfPpkd-k2Wrsb{margin-bottom:0;padding:0;border-bottom:0}.VfPpkd-Sx9Kwc-OWXEXe-n9oEIb.VfPpkd-Sx9Kwc-OWXEXe-s2gQvd .VfPpkd-k2Wrsb{border-bottom:0;margin-bottom:0}.VfPpkd-Sx9Kwc-OWXEXe-n9oEIb .VfPpkd-zMU9ub-suEOdc-sM5MNb{top:5px}.VfPpkd-Sx9Kwc-OWXEXe-n9oEIb.VfPpkd-Sx9Kwc-OWXEXe-s2gQvd .VfPpkd-T0kwCb{border-top:1px solid transparent}@media screen and (forced-colors:active){.VfPpkd-Sx9Kwc-OWXEXe-n9oEIb.VfPpkd-Sx9Kwc-OWXEXe-s2gQvd .VfPpkd-T0kwCb{border-top-color:CanvasText}}.VfPpkd-Sx9Kwc-OWXEXe-n9oEIb-OWXEXe-diJVc .VfPpkd-zMU9ub-suEOdc-sM5MNb{margin-top:4px}.VfPpkd-Sx9Kwc-OWXEXe-n9oEIb-OWXEXe-diJVc.VfPpkd-Sx9Kwc-OWXEXe-s2gQvd .VfPpkd-zMU9ub-suEOdc-sM5MNb{margin-top:0}.VfPpkd-cnG4Wd{-webkit-box-flex:1;-webkit-flex-grow:1;flex-grow:1;box-sizing:border-box;margin:0;overflow:auto}.VfPpkd-cnG4Wd>:first-child{margin-top:0}.VfPpkd-cnG4Wd>:last-child{margin-bottom:0}.VfPpkd-k2Wrsb+.VfPpkd-cnG4Wd,.VfPpkd-oclYLd+.VfPpkd-cnG4Wd{padding-top:0}.VfPpkd-Sx9Kwc-OWXEXe-s2gQvd .VfPpkd-k2Wrsb+.VfPpkd-cnG4Wd{padding-top:8px;padding-bottom:8px}.VfPpkd-cnG4Wd .VfPpkd-StrnGf-rymPhb:first-child:last-child{padding:6px 0 0}.VfPpkd-Sx9Kwc-OWXEXe-s2gQvd .VfPpkd-cnG4Wd .VfPpkd-StrnGf-rymPhb:first-child:last-child{padding:0}.VfPpkd-T0kwCb{display:-webkit-box;display:-webkit-flex;display:flex;position:relative;-webkit-flex-shrink:0;flex-shrink:0;-webkit-flex-wrap:wrap;flex-wrap:wrap;-webkit-box-align:center;-webkit-align-items:center;align-items:center;-webkit-box-pack:end;-webkit-justify-content:flex-end;justify-content:flex-end;box-sizing:border-box;min-height:52px;margin:0;padding:8px;border-top:1px solid transparent}@media screen and (forced-colors:active){.VfPpkd-T0kwCb{border-top-color:CanvasText}}.VfPpkd-Sx9Kwc-OWXEXe-eu7FSc .VfPpkd-T0kwCb{-webkit-box-orient:vertical;-webkit-box-direction:normal;-webkit-flex-direction:column;flex-direction:column;-webkit-box-align:end;-webkit-align-items:flex-end;align-items:flex-end}.VfPpkd-M1klYe{margin-left:8px;margin-right:0;max-width:100%;text-align:right}[dir=rtl] .VfPpkd-M1klYe,.VfPpkd-M1klYe[dir=rtl]{margin-left:0;margin-right:8px}.VfPpkd-M1klYe:first-child{margin-left:0;margin-right:0}[dir=rtl] .VfPpkd-M1klYe:first-child,.VfPpkd-M1klYe:first-child[dir=rtl]{margin-left:0;margin-right:0}[dir=rtl] .VfPpkd-M1klYe,.VfPpkd-M1klYe[dir=rtl]{text-align:left}.VfPpkd-Sx9Kwc-OWXEXe-eu7FSc .VfPpkd-M1klYe:not(:first-child){margin-top:12px}.VfPpkd-Sx9Kwc-OWXEXe-FNFY6c,.VfPpkd-Sx9Kwc-OWXEXe-uGFO6d,.VfPpkd-Sx9Kwc-OWXEXe-FnSee{display:-webkit-box;display:-webkit-flex;display:flex}.VfPpkd-Sx9Kwc-OWXEXe-uGFO6d .VfPpkd-IE5DDf{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.VfPpkd-Sx9Kwc-OWXEXe-uGFO6d .VfPpkd-wzTsW{-webkit-transition:opacity 75ms linear,-webkit-transform .15s 0ms cubic-bezier(0,0,.2,1);transition:opacity 75ms linear,-webkit-transform .15s 0ms cubic-bezier(0,0,.2,1);transition:opacity 75ms linear,transform .15s 0ms cubic-bezier(0,0,.2,1);transition:opacity 75ms linear,transform .15s 0ms cubic-bezier(0,0,.2,1),-webkit-transform .15s 0ms cubic-bezier(0,0,.2,1)}.VfPpkd-Sx9Kwc-OWXEXe-FnSee .VfPpkd-IE5DDf,.VfPpkd-Sx9Kwc-OWXEXe-FnSee .VfPpkd-wzTsW{-webkit-transition:opacity 75ms linear;transition:opacity 75ms linear}.VfPpkd-Sx9Kwc-OWXEXe-FnSee .VfPpkd-wzTsW,.VfPpkd-Sx9Kwc-OWXEXe-FnSee .VfPpkd-P5QLlc{-webkit-transform:none;transform:none}.VfPpkd-Sx9Kwc-OWXEXe-RTQbk .VfPpkd-IE5DDf{-webkit-transition:none;transition:none;opacity:1}.VfPpkd-Sx9Kwc-OWXEXe-FNFY6c .VfPpkd-IE5DDf,.VfPpkd-Sx9Kwc-OWXEXe-FNFY6c .VfPpkd-wzTsW{opacity:1}.VfPpkd-Sx9Kwc-OWXEXe-FNFY6c .VfPpkd-P5QLlc{-webkit-transform:none;transform:none}.VfPpkd-Sx9Kwc-OWXEXe-FNFY6c.VfPpkd-P5QLlc-GGAcbc-OWXEXe-TSZdd .VfPpkd-P5QLlc-GGAcbc{opacity:1}.VfPpkd-Sx9Kwc-OWXEXe-FNFY6c.VfPpkd-P5QLlc-GGAcbc-OWXEXe-wJB69c .VfPpkd-P5QLlc-GGAcbc{-webkit-transition:opacity 75ms linear;transition:opacity 75ms linear}.VfPpkd-Sx9Kwc-OWXEXe-FNFY6c.VfPpkd-P5QLlc-GGAcbc-OWXEXe-eo9XGd .VfPpkd-P5QLlc-GGAcbc{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.VfPpkd-P5QLlc-GGAcbc{display:none;opacity:0;position:absolute;width:100%;height:100%;z-index:1}.VfPpkd-P5QLlc-GGAcbc-OWXEXe-TSZdd .VfPpkd-P5QLlc-GGAcbc,.VfPpkd-P5QLlc-GGAcbc-OWXEXe-eo9XGd .VfPpkd-P5QLlc-GGAcbc,.VfPpkd-P5QLlc-GGAcbc-OWXEXe-wJB69c .VfPpkd-P5QLlc-GGAcbc{display:block}.VfPpkd-Sx9Kwc-XuHpsb-pGuBYc{overflow:hidden}.VfPpkd-Sx9Kwc-OWXEXe-di8rgd-bN97Pc-QFlW2 .VfPpkd-cnG4Wd{padding:0}.VfPpkd-Sx9Kwc-OWXEXe-vOE8Lb .VfPpkd-wzTsW .VfPpkd-zMU9ub-suEOdc-sM5MNb{right:12px;top:9px;position:absolute;z-index:1}.VfPpkd-IE5DDf-OWXEXe-uIDLbb{pointer-events:none}.VfPpkd-IE5DDf-OWXEXe-uIDLbb .VfPpkd-IE5DDf,.VfPpkd-IE5DDf-OWXEXe-uIDLbb .VfPpkd-P5QLlc-GGAcbc{display:none}.cC1eCc{z-index:2001}.cC1eCc .VfPpkd-k2Wrsb{color:#3c4043}.cC1eCc .VfPpkd-cnG4Wd{color:#5f6368}.cC1eCc .VfPpkd-zMU9ub{color:rgb(95,99,104)}.cC1eCc .VfPpkd-zMU9ub .VfPpkd-Bz112c-Jh9lGc::before,.cC1eCc .VfPpkd-zMU9ub .VfPpkd-Bz112c-Jh9lGc::after{background-color:rgb(95,99,104);background-color:var(--mdc-ripple-color,rgb(95,99,104))}.cC1eCc .VfPpkd-zMU9ub:hover .VfPpkd-Bz112c-Jh9lGc::before,.cC1eCc .VfPpkd-zMU9ub.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Bz112c-Jh9lGc::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.cC1eCc .VfPpkd-zMU9ub.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Bz112c-Jh9lGc::before,.cC1eCc .VfPpkd-zMU9ub:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Bz112c-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.cC1eCc .VfPpkd-zMU9ub:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Bz112c-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.cC1eCc .VfPpkd-zMU9ub:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Bz112c-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-press-opacity,.12)}.cC1eCc .VfPpkd-zMU9ub.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.12)}.cC1eCc .VfPpkd-IE5DDf,.cC1eCc .VfPpkd-P5QLlc-GGAcbc{background-color:rgba(32,33,36,.6)}.cC1eCc .VfPpkd-P5QLlc{background-color:#fff}.cC1eCc .VfPpkd-P5QLlc{border-width:0;box-shadow:0 1px 3px 0 rgba(60,64,67,.3),0 4px 8px 3px rgba(60,64,67,.15)}.cC1eCc .VfPpkd-P5QLlc .VfPpkd-BFbNVe-bF1uUb{opacity:0}.cC1eCc .VfPpkd-P5QLlc{border-radius:8px}.cC1eCc .VfPpkd-T0kwCb{padding-top:2px;padding-bottom:2px}.cC1eCc .VfPpkd-T0kwCb .VfPpkd-RLmnJb{top:-6px;-webkit-transform:none;transform:none}.cC1eCc .VfPpkd-k2Wrsb{font-family:"Google Sans",Roboto,Arial,sans-serif;line-height:1.5rem;font-size:1rem;letter-spacing:.00625em;font-weight:500;padding-bottom:13px}.cC1eCc .VfPpkd-cnG4Wd{font-family:Roboto,Arial,sans-serif;line-height:1.25rem;font-size:.875rem;letter-spacing:.0142857143em;font-weight:400}.cC1eCc .VfPpkd-T0kwCb .VfPpkd-LgbsSe+.VfPpkd-LgbsSe{margin-left:8px}.cC1eCc.VfPpkd-Sx9Kwc-OWXEXe-n9oEIb .VfPpkd-k2Wrsb{font-family:"Google Sans",Roboto,Arial,sans-serif;line-height:1.5rem;font-size:1.125rem;letter-spacing:0;font-weight:400;padding-bottom:0}.iGu0Be{text-align:center}[dir=rtl] .iGu0Be,.iGu0Be[dir=rtl]{text-align:center}.nE3Lu{color:rgb(26,115,232);height:24px;width:24px}.nE3Lu::after{content:"";display:block}.bYmtV .VfPpkd-P5QLlc{background-color:#fff;color:rgb(95,99,104);font-family:roboto,"Noto Sans Myanmar UI",arial,sans-serif;letter-spacing:0.25px}.bYmtV .VfPpkd-k2Wrsb{color:rgb(32,33,36);font-family:"Google Sans","Noto Sans Myanmar UI",arial,sans-serif;font-size:20px;font-weight:500;letter-spacing:0.25px;line-height:1.3333}.bYmtV .VfPpkd-cnG4Wd{font-family:roboto,"Noto Sans Myanmar UI",arial,sans-serif;font-size:14px;letter-spacing:0.25px;line-height:1.4286;padding-bottom:0}.bYmtV .VfPpkd-T0kwCb{padding:0 24px 8px 24px}.bYmtV .VfPpkd-Bz112c-LgbsSe .VfPpkd-Bz112c-Jh9lGc::before,.bYmtV .VfPpkd-Bz112c-LgbsSe .VfPpkd-Bz112c-Jh9lGc::after{border-radius:4px}.bYmtV.Zttm2{border-radius:0}.bYmtV.Zttm2 .VfPpkd-P5QLlc{height:100vh;max-height:none;max-width:none;width:100vw}.bYmtV.Zttm2 .AH8Npc{height:100%;width:100%}.bYmtV .CJRWze{color:rgb(95,99,104);font-family:roboto,"Noto Sans Myanmar UI",arial,sans-serif;-webkit-box-flex:1;-webkit-flex-grow:1;flex-grow:1;font-size:12px;font-weight:400;padding-left:16px}.CwHtnf{border:none;color-scheme:normal;display:block;height:100%;padding:0;width:100%}.bYmtV .CxRgyd{margin-left:0;margin-right:0;padding-left:0;padding-right:0}:root{--wf-color-warning-bg:#fff0d1;--wf-color-warning-icon:#f09d00;--wf-color-warning-text:#421f00}@media screen and (prefers-color-scheme:dark){:root{--wf-color-warning-bg:#754200;--wf-color-warning-icon:#ffdf99;--wf-color-warning-text:#fff0d1}}.NAHnJe:not(:first-child){margin-top:8px}.NAHnJe:not(:last-child){margin-bottom:8px}.wClb9e{color:var(--gm3-sys-color-on-surface,#1f1f1f);margin-bottom:8px;font-family:Google Sans,Roboto,Noto Sans Myanmar UI,Arial,sans-serif;font-weight:400;font-size:1rem;letter-spacing:0rem;line-height:1.5rem}.XQGu9e{padding-bottom:16px;padding-left:16px;padding-right:16px}.eoX0T{width:100%}.eoX0T.MyuJQe{margin-bottom:8px;border-top-left-radius:20px;border-top-right-radius:20px;border-bottom-left-radius:20px;border-bottom-right-radius:20px}.gTwoD{-webkit-box-align:start;-webkit-align-items:flex-start;align-items:flex-start;display:-webkit-inline-box;display:-webkit-inline-flex;display:inline-flex;-webkit-box-pack:justify;-webkit-justify-content:space-between;justify-content:space-between;padding:0;width:100%}.lWCUk{background-color:var(--gm3-sys-color-surface-container,#f0f4f9);border-radius:4px;margin:2px 0;-webkit-transition:border-radius .1s cubic-bezier(.2,0,0,1);transition:border-radius .1s cubic-bezier(.2,0,0,1)}.lWCUk:first-child{margin-top:0;border-top-left-radius:20px;border-top-right-radius:20px}.lWCUk:last-child{margin-bottom:0;border-bottom-left-radius:20px;border-bottom-right-radius:20px}.lWCUk .lWCUk{background:var(--gm3-sys-color-surface-bright,#fff);border-radius:4px}.lWCUk .lWCUk:first-child{border-top-left-radius:16px;border-top-right-radius:16px}.lWCUk .lWCUk:last-child{border-bottom-left-radius:16px;border-bottom-right-radius:16px}.lWCUk.KKjvXb:not(.RDPZE){border-radius:28px}.lWCUk>.gTwoD{padding-left:16px;padding-right:16px}.lWCUk>.gTwoD.NEk0Ve{padding-left:8px}.lWCUk>.gTwoD.zVkt0c{padding-left:4px}.lWCUk>.gTwoD.NEk0Ve.kS4AXe{padding-left:16px;padding-right:8px}.lWCUk>.gTwoD.zVkt0c.kS4AXe{padding-left:16px;padding-right:4px}.lWCUk>.gTwoD:has(.GnLI0e.o96OHc){padding-left:0}.GnLI0e{cursor:pointer;display:-webkit-box;display:-webkit-flex;display:flex;-webkit-box-flex:1;-webkit-flex-grow:1;flex-grow:1;padding:18px 0}.gTwoD.NEk0Ve .GnLI0e{margin-left:8px}.gTwoD.zVkt0c .GnLI0e{margin-left:4px}.gTwoD.kS4AXe .GnLI0e{margin-left:0}.GnLI0e:has(.sQ1LEb){padding-bottom:12px;padding-top:12px}.GnLI0e,.GnLI0e .XZVJqc{min-width:0;width:100%}.GnLI0e .XZVJqc{display:inline-block;-webkit-box-flex:1;-webkit-flex-grow:1;flex-grow:1;text-align:left}.GnLI0e .kM29Gb{color:var(--gm3-sys-color-on-surface,#1f1f1f);font-family:Google Sans,Roboto,Noto Sans Myanmar UI,Arial,sans-serif;font-size:1rem;font-weight:400;letter-spacing:0rem;line-height:1.5rem}.GnLI0e .sQ1LEb{color:var(--gm3-sys-color-on-surface-variant,#444746);font-family:Google Sans,Roboto,Noto Sans Myanmar UI,Arial,sans-serif;font-size:0.875rem;font-weight:400;letter-spacing:0rem;line-height:1.25rem}.GnLI0e .kM29Gb,.GnLI0e .sQ1LEb{display:block;overflow:hidden;text-overflow:ellipsis;width:100%}.eoX0T.RDPZE>.gTwoD .GnLI0e:not(.o96OHc){cursor:default;opacity:0.38}.GnLI0e.o96OHc{background:transparent;border:0;color:inherit;-webkit-box-pack:justify;-webkit-justify-content:space-between;justify-content:space-between;text-decoration:none;--gm3-focus-ring-outward-target-shape-start-start:4px;--gm3-focus-ring-outward-target-shape-start-end:4px;--gm3-focus-ring-outward-target-shape-end-end:4px;--gm3-focus-ring-outward-target-shape-end-start:4px}.GnLI0e.o96OHc{position:relative}.GnLI0e.o96OHc::before{background:var(--gm3-sys-color-on-surface,#1f1f1f);content:"";opacity:0;position:absolute;pointer-events:none}.GnLI0e.o96OHc:hover::before{opacity:0.08}.GnLI0e.o96OHc:focus:not(:hover)::before,.GnLI0e.o96OHc.u3bW4e::before{opacity:0.1}.GnLI0e.o96OHc:active::before,.GnLI0e.o96OHc.qs41qe::before{opacity:0.1}.GnLI0e.o96OHc::before{border-radius:4px;height:100%;left:-16px;right:0;top:0}.GnLI0e.o96OHc:focus:not(:hover)::before,.GnLI0e.o96OHc.u3bW4e::before{display:none}.GnLI0e.o96OHc:focus-visible{outline:none;--gm3-focus-ring-outward-display:block}.lWCUk .GnLI0e.o96OHc{padding-left:16px}.lWCUk .GnLI0e.o96OHc::before{left:0}.GnLI0e.o96OHc:has(.sQ1LEb){padding-bottom:12px;padding-top:12px}.eoX0T:first-of-type .GnLI0e.o96OHc{--gm3-focus-ring-outward-target-shape-start-start:20px}.eoX0T:first-of-type .GnLI0e.o96OHc::before{border-top-left-radius:20px}.eoX0T:last-of-type .GnLI0e.o96OHc{--gm3-focus-ring-outward-target-shape-end-start:20px}.eoX0T:last-of-type .GnLI0e.o96OHc::before{border-bottom-left-radius:20px}.lWCUk.KKjvXb .GnLI0e.o96OHc{--gm3-focus-ring-outward-target-shape-start-start:28px;--gm3-focus-ring-outward-target-shape-end-start:28px}.lWCUk.KKjvXb .GnLI0e.o96OHc::before{border-top-left-radius:28px;border-bottom-left-radius:28px}.GnLI0e.o96OHc::after{background:var(--gm3-sys-color-outline,#747775);content:"";display:block;height:40px;position:absolute;right:0;top:11px;width:1px}.gTwoD.NEk0Ve .GnLI0e.o96OHc{margin-right:8px}.gTwoD.zVkt0c .GnLI0e.o96OHc{margin-right:4px}.GnLI0e:has(.sQ1LEb).o96OHc::after{position:relative;top:calc(1.375rem - 20px)}.UjRYsb{color:var(--gm3-sys-color-on-surface-variant,#444746);min-height:24px;min-width:24px;position:relative;top:-1px}.eoX0T .UjRYsb{margin-left:16px}.gTwoD.kS4AXe .UjRYsb{margin-left:0;margin-right:16px}.uxn3Pd{fill:var(--gm3-sys-color-on-surface,#1f1f1f);margin-right:16px;min-height:24px;min-width:24px;position:relative}.GnLI0e:has(.sQ1LEb)>.UjRYsb,.GnLI0e:has(.sQ1LEb)>.uxn3Pd{position:relative;top:calc((2.75rem - 24px)/2)}.xCCdfe{position:relative}.xCCdfe.NEk0Ve{top:calc(18px - ((40px - 1.5rem)/2))}.xCCdfe.zVkt0c{top:calc(18px - ((48px - 1.5rem)/2))}.xCCdfe.Msforc{padding-left:16px;top:calc(18px - ((32px - 1.5rem)/2));--gm3-sys-color-on-surface-rgb:31,31,31}@media screen and (prefers-color-scheme:dark){.xCCdfe.Msforc{--gm3-sys-color-on-surface-rgb:227,227,227}}.gTwoD:has(.sQ1LEb) .xCCdfe.NEk0Ve{position:relative;top:calc(1.375rem - 10px)}.gTwoD:has(.sQ1LEb) .xCCdfe.zVkt0c{position:relative;top:calc(1.375rem - 12px)}.gTwoD:has(.sQ1LEb) .xCCdfe.Msforc{padding-top:12px;position:relative;top:calc(1.375rem - 16px)}.A2WLNb{background:var(--gm3-sys-color-surface-container,#f0f4f9);border-radius:28px;margin:8px 0;-webkit-transition:border-radius .1s cubic-bezier(.2,0,0,1);transition:border-radius .1s cubic-bezier(.2,0,0,1)}.A2WLNb.jVwmLb{border-radius:20px;padding-bottom:0}.A2WLNb .WKpdi{-webkit-box-flex:1;-webkit-flex-grow:1;flex-grow:1}.A2WLNb .lWCUk{background:var(--gm3-sys-color-surface-bright,#fff);border-radius:4px}.A2WLNb .lWCUk:first-child{border-top-left-radius:16px;border-top-right-radius:16px}.A2WLNb .lWCUk:last-child{border-bottom-left-radius:16px;border-bottom-right-radius:16px}.A2WLNb .lWCUk.KKjvXb:not(.RDPZE){border-radius:28px}.KrF7fd{-webkit-box-align:start;-webkit-align-items:flex-start;align-items:flex-start;background:transparent;border:0;display:-webkit-inline-box;display:-webkit-inline-flex;display:inline-flex;-webkit-box-pack:justify;-webkit-justify-content:space-between;justify-content:space-between;padding-left:16px;padding-right:16px;width:100%;text-decoration:none;--gm3-focus-ring-outward-target-shape-start-start:28px;--gm3-focus-ring-outward-target-shape-start-end:28px;--gm3-focus-ring-outward-target-shape-end-end:28px;--gm3-focus-ring-outward-target-shape-end-start:28px}.KrF7fd{position:relative}.KrF7fd::before{background:var(--gm3-sys-color-on-surface,#1f1f1f);content:"";opacity:0;position:absolute;pointer-events:none}.KrF7fd:hover::before{opacity:0.08}.KrF7fd:focus:not(:hover)::before,.KrF7fd.u3bW4e::before{opacity:0.1}.KrF7fd:active::before,.KrF7fd.qs41qe::before{opacity:0.1}.KrF7fd::before{border-radius:28px;height:100%;left:0;right:0;top:0}.KrF7fd:focus:not(:hover)::before,.KrF7fd.u3bW4e::before{display:none}.KrF7fd:focus-visible{outline:none;--gm3-focus-ring-outward-display:block}.A2WLNb.jVwmLb .KrF7fd::before{border-radius:20px}.KrF7fd .RwGqvd{margin-left:0;margin-right:16px}.A2WLNb:has(.sQ1LEb) .RwGqvd{position:relative;top:calc((2.75rem - 24px)/2)}.A2WLNb .xIgdGc{-webkit-box-align:center;-webkit-align-items:center;align-items:center;background:var(--gm3-sys-color-secondary-container,#c2e7ff);border-radius:12px;display:-webkit-box;display:-webkit-flex;display:flex;height:24px;-webkit-box-pack:center;-webkit-justify-content:center;justify-content:center;min-width:24px}.A2WLNb.jVwmLb .xIgdGc{background:var(--gm3-sys-color-surface-bright,#fff)}.A2WLNb:has(.sQ1LEb) .xIgdGc{position:relative;top:calc((2.75rem - 24px)/2)}.A2WLNb .eZIgdb{fill:var(--gm3-sys-color-on-secondary-container,#004a77);-webkit-transform:rotate(180deg);transform:rotate(180deg)}.A2WLNb.jVwmLb .eZIgdb{fill:var(--gm3-sys-color-on-surface-variant,#444746);-webkit-transform:rotate(0);transform:rotate(0)}.jzGg7c{padding-bottom:16px;padding-left:16px;padding-right:16px}.A2WLNb.jVwmLb .jzGg7c{display:none}:root{--wf-tfs:calc(var(--c-tfs,32)/16*1rem);--wf-tfs-bp2:calc(var(--c-tfs,36)/16*1rem);--wf-tfs-bp3:calc(var(--c-tfs,36)/16*1rem);--wf-tfs-bp5:calc(var(--c-tfs,44)/16*1rem);--wf-stfs:calc(var(--c-stfs,16)/16*1rem);--wf-stfs-bp5:calc(var(--c-stfs,16)/16*1rem)}.B6L7ke{height:25vh;margin:auto -24px;min-height:110px;padding-left:24px;padding-right:24px;position:relative}.SCAiR{height:25vh;margin:auto -24px;min-height:110px;padding-left:24px;padding-right:24px;position:relative;overflow:hidden}.JtUbMb,.Nny6ue{display:block;height:100%;margin:0 auto;object-fit:contain;width:100%}@media (min-width:450px){.B6L7ke{margin:auto -40px;padding-left:40px;padding-right:40px}}@media (min-width:601px){.B6L7ke{height:150px}}.B6L7ke.Irjbwb{height:auto}.B6L7ke.IiQozc{text-align:center}.xh7Wmd{height:25vh;max-width:100%;min-height:110px;position:relative;-webkit-transform:translate(-43%,-3%);transform:translate(-43%,-3%);z-index:3}@media (min-width:601px){.xh7Wmd{height:150px}}.B6L7ke.FnDdB{height:auto}.B6L7ke.FnDdB .xh7Wmd{height:auto;max-width:312px;width:100%}.B6L7ke.FnDdB.zpCp3 .xh7Wmd{max-width:unset}.B6L7ke.IiQozc .xh7Wmd{-webkit-transform:none;transform:none}.B6L7ke.aJJFde .xh7Wmd{left:-100%;margin:auto;position:absolute;right:-100%;-webkit-transform:translate(0,-3%);transform:translate(0,-3%)}.B6L7ke.Irjbwb .xh7Wmd{height:auto;width:100%}.p17Urb{background-image:-webkit-linear-gradient(to bottom,rgba(233,233,233,0) 0%,rgba(233,233,233,0) 62.22%,rgba(233,233,233,1) 40.22%,rgba(233,233,233,0) 100%);background-image:linear-gradient(to bottom,rgba(233,233,233,0) 0%,rgba(233,233,233,0) 62.22%,rgba(233,233,233,1) 40.22%,rgba(233,233,233,0) 100%);height:100%;left:0;overflow:hidden;position:absolute;right:0;top:0;z-index:2}.p17Urb::after,.p17Urb::before{content:"";display:block;height:100%;min-width:110px;position:absolute;right:-10%;-webkit-transform:rotate(-104deg);transform:rotate(-104deg);width:25vh;z-index:2}@media (min-width:601px){.p17Urb::after,.p17Urb::before{width:150px}}.p17Urb::before{background-image:-webkit-linear-gradient(to bottom,rgba(243,243,243,0) 0%,rgba(243,243,243,.9) 100%);background-image:linear-gradient(to bottom,rgba(243,243,243,0) 0%,rgba(243,243,243,.9) 100%);bottom:-10%}.p17Urb::after{background-image:-webkit-linear-gradient(to bottom,rgba(255,255,255,0) 0%,rgba(255,255,255,.9) 100%);background-image:linear-gradient(to bottom,rgba(255,255,255,0) 0%,rgba(255,255,255,.9) 100%);bottom:-80%}.DrceJe{height:auto}.yb5i2e{-webkit-transform:translate(-9%,-3%);transform:translate(-9%,-3%)}.hNLjwb{-webkit-transform:translate(9%,-3%);transform:translate(9%,-3%)}.ulNYne{left:-40%;margin:auto;max-height:230px;position:absolute;right:0;top:-3%;-webkit-transform:none;transform:none}.F8EZte{-webkit-transform:translate(24px,0);transform:translate(24px,0)}.eMXECe{-webkit-transform:translate(0,0);transform:translate(0,0)}.B6L7ke.i1L7v{height:15vh;max-height:137px;min-height:112px;padding-bottom:12px}.B6L7ke.i1L7v .xh7Wmd{max-height:100%;min-height:100%}.B6L7ke.j1zy9{height:auto}.B6L7ke.j1zy9 .xh7Wmd{height:auto;max-width:432px}.PeAiAb{max-width:300px}.MWnvBb.WS4XDd{border:0;max-height:1rem;padding:0 2px;vertical-align:middle;width:auto}.IqauWe{border:0;object-fit:contain}.IqauWe.WS4XDd{border:0;max-height:1rem;padding:0 2px;vertical-align:middle;width:auto}.q4Wquf,.nfoC7c{display:block;height:25vh;position:relative}@media (min-width:600px){.q4Wquf,.nfoC7c{height:150px}}.q4Wquf.Irjbwb{height:auto}@media screen and (prefers-color-scheme:dark){.q4Wquf:not(.GtvzYd){display:none}}.nfoC7c{margin:0;overflow:hidden}.PwpMUe,.lVUmD{display:block;height:100%;margin:0 auto;object-fit:contain;width:100%}.St9mde{display:block;height:100%;max-width:100%;min-height:110px;position:relative;-webkit-transform:translate(-43%,-3%);transform:translate(-43%,-3%);width:auto;z-index:3}.wsArZ[data-ss-mode="1"] .q4Wquf,.wsArZ[data-ss-mode="1"] .St9mde{height:auto;width:100%}.wsArZ[data-ss-mode="1"] .St9mde{max-width:400px}@media (min-width:600px) and (orientation:landscape),all and (min-width:1600px){.NQ5OL .q4Wquf,.NQ5OL .St9mde{height:auto;width:100%}.NQ5OL .St9mde{max-width:400px}}.q4Wquf.NWba7e,.q4Wquf.NWba7e .St9mde{height:auto}.q4Wquf.NWba7e .St9mde{height:auto;max-width:312px;width:100%}.q4Wquf.NWba7e.zpCp3 .St9mde{max-width:unset}.q4Wquf.IiQozc .St9mde{margin:0 auto;-webkit-transform:none;transform:none}.q4Wquf.Irjbwb .St9mde{height:auto;width:100%}.q4Wquf.EEeaqf .St9mde{max-height:144px;max-width:144px}.SnAaEd{background-image:-webkit-gradient(linear,left top,left bottom,from(rgba(233,233,233,0)),color-stop(62.22%,rgba(233,233,233,0)),color-stop(40.22%,rgb(233,233,233)),to(rgba(233,233,233,0)));background-image:-webkit-linear-gradient(top,rgba(233,233,233,0) 0,rgba(233,233,233,0) 62.22%,rgb(233,233,233) 40.22%,rgba(233,233,233,0) 100%);background-image:linear-gradient(to bottom,rgba(233,233,233,0) 0,rgba(233,233,233,0) 62.22%,rgb(233,233,233) 40.22%,rgba(233,233,233,0) 100%);height:100%;left:0;overflow:hidden;position:absolute;right:0;top:0;z-index:2}@media screen and (prefers-color-scheme:dark){.SnAaEd{display:none}}.SnAaEd::after,.SnAaEd::before{content:"";display:block;height:100%;min-width:110px;position:absolute;right:-10%;-webkit-transform:rotate(-104deg);transform:rotate(-104deg);width:25vh;z-index:2}@media (min-width:600px){.SnAaEd::after,.SnAaEd::before{width:150px}}.SnAaEd::before{background-image:-webkit-gradient(linear,left top,left bottom,from(rgba(243,243,243,0)),to(rgba(243,243,243,.9)));background-image:-webkit-linear-gradient(top,rgba(243,243,243,0) 0,rgba(243,243,243,.9) 100%);background-image:linear-gradient(to bottom,rgba(243,243,243,0) 0,rgba(243,243,243,.9) 100%);bottom:-10%}.SnAaEd::after{background-image:-webkit-gradient(linear,left top,left bottom,from(rgba(255,255,255,0)),to(rgba(255,255,255,.9)));background-image:-webkit-linear-gradient(top,rgba(255,255,255,0) 0,rgba(255,255,255,.9) 100%);background-image:linear-gradient(to bottom,rgba(255,255,255,0) 0,rgba(255,255,255,.9) 100%);bottom:-80%}.wsArZ[data-ss-mode="1"] .SnAaEd~.St9mde{width:auto}@media (min-width:600px) and (orientation:landscape),all and (min-width:1600px){.NQ5OL .SnAaEd~.St9mde{width:auto}}.RHNWk .St9mde{height:auto}@media (min-width:600px) and (orientation:landscape),all and (min-width:1600px){.NQ5OL .RHNWk .St9mde{width:115px}}.cf660d .St9mde{-webkit-transform:translate(-9%,-3%);transform:translate(-9%,-3%)}.tUhwwc .St9mde{margin:auto;max-height:230px;right:0;top:-3%;-webkit-transform:none;transform:none}.Jkvqxd .St9mde{-webkit-transform:translate(9%,-3%);transform:translate(9%,-3%)}.onc8Ic .St9mde{-webkit-transform:translate(var(
    --c-ps-s,24px
  ),0);transform:translate(var(
    --c-ps-s,24px
  ),0)}.WA89Yb .St9mde{-webkit-transform:translate(0,0);transform:translate(0,0)}.wsArZ[data-ss-mode="1"] .XEN8Yb .St9mde{max-width:115px}@media (min-width:600px) and (orientation:landscape),all and (min-width:1600px){.NQ5OL .XEN8Yb .St9mde{max-width:115px}}.IsSr6b .St9mde{max-width:300px}.mmskdd .St9mde{-webkit-transform:none;transform:none}.Qk3oof.WS4XDd{border:0;max-height:1.4285714286em;padding:0 2px;vertical-align:middle;width:auto}.uHLU0{border:0;object-fit:contain}.uHLU0.WS4XDd{border:0;max-height:1.4285714286em;padding:0 2px;vertical-align:middle;width:auto}.Dzz9Db,.GpMPBe{display:block;height:25vh;position:relative}@media (min-width:600px){.Dzz9Db,.GpMPBe{height:150px}}@media screen and (prefers-color-scheme:dark){.Dzz9Db:not(.GtvzYd){display:none}}.Dzz9Db.Irjbwb{height:auto}.GpMPBe{margin:0;overflow:hidden}.UFQPDd,.JNOvdd{display:block;height:100%;margin:0 auto;object-fit:contain;width:100%}.f4ZpM{display:block;height:100%;max-width:100%;min-height:110px;position:relative;-webkit-transform:translate(-43%,-3%);transform:translate(-43%,-3%);width:auto;z-index:3}.wsArZ[data-ss-mode="1"] .Dzz9Db,.wsArZ[data-ss-mode="1"] .f4ZpM{height:auto;width:100%}.wsArZ[data-ss-mode="1"] .f4ZpM{max-width:400px}@media (min-width:600px) and (orientation:landscape),all and (min-width:1600px){.NQ5OL .Dzz9Db,.NQ5OL .f4ZpM{height:auto;width:100%}.NQ5OL .f4ZpM{max-width:400px}}.Dzz9Db.utFBGf,.Dzz9Db.utFBGf .f4ZpM{height:auto}.Dzz9Db.utFBGf .f4ZpM{height:auto;max-width:312px;width:100%}.Dzz9Db.utFBGf.zpCp3 .f4ZpM{max-width:unset}.Dzz9Db.IiQozc .f4ZpM{margin:0 auto;-webkit-transform:none;transform:none}.Dzz9Db.Irjbwb .f4ZpM{height:auto;width:100%}.Dzz9Db.EEeaqf .f4ZpM{max-height:144px;max-width:144px}.nPt1pc{background-image:-webkit-gradient(linear,left top,left bottom,from(rgba(233,233,233,0)),color-stop(62.22%,rgba(233,233,233,0)),color-stop(40.22%,rgb(233,233,233)),to(rgba(233,233,233,0)));background-image:-webkit-linear-gradient(top,rgba(233,233,233,0) 0,rgba(233,233,233,0) 62.22%,rgb(233,233,233) 40.22%,rgba(233,233,233,0) 100%);background-image:linear-gradient(to bottom,rgba(233,233,233,0) 0,rgba(233,233,233,0) 62.22%,rgb(233,233,233) 40.22%,rgba(233,233,233,0) 100%);height:100%;left:0;overflow:hidden;position:absolute;right:0;top:0;z-index:2}@media screen and (prefers-color-scheme:dark){.nPt1pc{display:none}}.nPt1pc::after,.nPt1pc::before{content:"";display:block;height:100%;min-width:110px;position:absolute;right:-10%;-webkit-transform:rotate(-104deg);transform:rotate(-104deg);width:25vh;z-index:2}@media (min-width:600px){.nPt1pc::after,.nPt1pc::before{width:150px}}.nPt1pc::before{background-image:-webkit-gradient(linear,left top,left bottom,from(rgba(243,243,243,0)),to(rgba(243,243,243,.9)));background-image:-webkit-linear-gradient(top,rgba(243,243,243,0) 0,rgba(243,243,243,.9) 100%);background-image:linear-gradient(to bottom,rgba(243,243,243,0) 0,rgba(243,243,243,.9) 100%);bottom:-10%}.nPt1pc::after{background-image:-webkit-gradient(linear,left top,left bottom,from(rgba(255,255,255,0)),to(rgba(255,255,255,.9)));background-image:-webkit-linear-gradient(top,rgba(255,255,255,0) 0,rgba(255,255,255,.9) 100%);background-image:linear-gradient(to bottom,rgba(255,255,255,0) 0,rgba(255,255,255,.9) 100%);bottom:-80%}.wsArZ[data-ss-mode="1"] .nPt1pc~.f4ZpM{width:auto}@media (min-width:600px) and (orientation:landscape),all and (min-width:1600px){.NQ5OL .nPt1pc~.f4ZpM{width:auto}}.ZS7CGc .f4ZpM{height:auto}@media (min-width:600px) and (orientation:landscape),all and (min-width:1600px){.NQ5OL .ZS7CGc .f4ZpM{width:115px}}.qiRZ5e .f4ZpM{-webkit-transform:translate(-9%,-3%);transform:translate(-9%,-3%)}.vIv7Gf .f4ZpM{margin:auto;max-height:230px;right:0;top:-3%;-webkit-transform:none;transform:none}.nvYXVd .f4ZpM{-webkit-transform:translate(9%,-3%);transform:translate(9%,-3%)}.uOhnzd .f4ZpM{-webkit-transform:translate(24px,0);transform:translate(24px,0)}.MsYMaf .f4ZpM{-webkit-transform:translate(0,0);transform:translate(0,0)}.wsArZ[data-ss-mode="1"] .YIi9qf .f4ZpM{max-width:115px}@media (min-width:600px) and (orientation:landscape),all and (min-width:1600px){.NQ5OL .YIi9qf .f4ZpM{max-width:115px}}.QG3Xbe .f4ZpM{max-width:300px}.F6gtje .f4ZpM{-webkit-transform:none;transform:none}.iHd3uf{display:-webkit-inline-box;display:-webkit-inline-flex;display:inline-flex}.iHd3uf.eLNT1d{display:none}.ceOhk{--gm3-button-filled-container-height:40px;--gm3-button-filled-container-shape:20px;--gm3-button-filled-label-text-weight:var(--c-afwt,500)}.WyRBD{--gm3-button-outlined-container-height:40px;--gm3-button-outlined-label-text-weight:var(--c-afwt,500);--gm3-button-outlined-container-shape:20px}.Xq56fd{--gm3-button-text-container-height:40px;--gm3-button-text-container-shape:20px;--gm3-button-text-label-text-weight:var(--c-afwt,500)}.hy0HVb{--gm3-button-filled-tonal-container-height:40px;--gm3-button-filled-tonal-container-shape:20px;--gm3-button-filled-tonal-label-text-weight:var(--c-afwt,500)}.ySLakb{margin:16px 0;outline:none}.ZfdVuf{margin:0 0}.ySLakb+.ySLakb:not(.ZfdVuf){margin-top:24px}.xe7Heb{margin-bottom:24px;margin-top:8px}.ySLakb:first-child{margin-top:0}.ySLakb:last-child{margin-bottom:0}.xHr6Xe{-webkit-box-align:center;-webkit-align-items:center;align-items:center;color:var(--gm3-sys-color-on-surface,#1f1f1f);display:-webkit-box;display:-webkit-flex;display:flex;margin-top:0;margin-bottom:0;padding:0 0 8px;font-family:Google Sans,Roboto,Noto Sans Myanmar UI,Arial,sans-serif;font-weight:400;font-size:1.25rem;letter-spacing:0rem;line-height:1.5rem}.xe7Heb>.Y9aYob .xHr6Xe{padding-bottom:12px}.ySLakb .xHr6Xe:has(.M0cpdd:empty),.i3HiPd.YFdWic .xHr6Xe,.Ci1RI .xHr6Xe{padding-bottom:0}.i3HiPd{border-radius:8px;padding:16px}.i3HiPd>:first-child{margin-top:0}.i3HiPd>:last-child{margin-bottom:0}.i3HiPd>.Y9aYob .xHr6Xe{font-family:Google Sans,Roboto,Noto Sans Myanmar UI,Arial,sans-serif;font-weight:500;font-size:1rem;letter-spacing:0rem;line-height:1.5rem}.i3HiPd.sj692e .xHr6Xe,.i3HiPd.sj692e .F4tG3e{color:var(--gm3-sys-color-on-primary-container,#0842a0)}.i3HiPd.Xq8bDe .xHr6Xe,.i3HiPd.Xq8bDe .F4tG3e{color:var(--gm3-sys-color-on-error-container,#8c1d18)}.i3HiPd.rNe0id .xHr6Xe,.i3HiPd.rNe0id .F4tG3e{color:var(
    --wf-color-warning-text,#421f00
  )}.i3HiPd.YFdWic .Y9aYob,.i3HiPd.YFdWic .F4tG3e{margin-left:64px;width:calc(100% - 48px - 16px)}.i3HiPd.YFdWic .F4tG3e{color:var(--gm3-sys-color-on-surface-variant,#444746)}.i3HiPd.YFdWic .xHr6Xe{color:var(--gm3-sys-color-on-surface,#1f1f1f)}.i3HiPd.YFdWic:not(.S7S4N) .Y9aYob{margin-left:0;width:0}.i3HiPd.sj692e{background:var(--gm3-sys-color-primary-container,#d3e3fd)}.i3HiPd.Xq8bDe{background:var(--gm3-sys-color-error-container,#f9dedc)}.i3HiPd.rNe0id{background:var(
    --wf-color-warning-bg,#fff0d1
  )}.i3HiPd.YFdWic{background:var(--gm3-sys-color-surface-container-low,#f8fafd);min-height:80px;position:relative}.i3HiPd:not(.S7S4N){display:-webkit-box;display:-webkit-flex;display:flex}.ySLakb.eLNT1d{display:none}.Ci1RI{background:var(--gm3-sys-color-surface-container,#f0f4f9);border-radius:20px;padding:16px}.Ci1RI>.Y9aYob .xHr6Xe{color:var(--gm3-sys-color-on-surface,#1f1f1f)}.Ci1RI .Zy76pd .snByac,.Ci1RI .Zy76pd.u3bW4e .snByac{background-color:var(--gm3-sys-color-surface-container,#f0f4f9)}.Ci1RI .rcBv3{display:-webkit-box;display:-webkit-flex;display:flex;-webkit-box-pack:end;-webkit-justify-content:flex-end;justify-content:flex-end;margin-top:16px}.Ci1RI .rcBv3 .hy0HVb{margin-bottom:0;margin-top:0;--gm3-button-filled-tonal-leading-space:16px;--gm3-button-filled-tonal-trailing-space:16px}.Ci1RI .F4tG3e .lWCUk{background:var(--gm3-sys-color-surface-bright,#fff);border-radius:4px}.Ci1RI .F4tG3e .lWCUk:first-child{border-top-left-radius:16px;border-top-right-radius:16px}.Ci1RI .F4tG3e .lWCUk:last-child{border-bottom-left-radius:16px;border-bottom-right-radius:16px}.ZfdVuf{border-bottom:1px solid var(--gm3-sys-color-outline-variant,#c4c7c5);display:-webkit-box;display:-webkit-flex;display:flex;-webkit-box-orient:vertical;-webkit-box-direction:normal;-webkit-flex-direction:column;flex-direction:column}.ZfdVuf .ZfdVuf:last-child{border-bottom:0}.ZfdVuf .Y9aYob{cursor:pointer;--gm3-focus-ring-outward-target-shape-start-start:8px;--gm3-focus-ring-outward-target-shape-start-end:8px;--gm3-focus-ring-outward-target-shape-end-end:8px;--gm3-focus-ring-outward-target-shape-end-start:8px}.ZfdVuf .Y9aYob{position:relative}.ZfdVuf .Y9aYob::before{background:var(--gm3-sys-color-on-surface,#1f1f1f);content:"";opacity:0;position:absolute;pointer-events:none}.ZfdVuf .Y9aYob:hover::before{opacity:0.08}.ZfdVuf .Y9aYob:focus:not(:hover)::before,.ZfdVuf .Y9aYob.u3bW4e::before{opacity:0.1}.ZfdVuf .Y9aYob:active::before,.ZfdVuf .Y9aYob.qs41qe::before{opacity:0.1}.ZfdVuf .Y9aYob::before{border-radius:8px;inset:0 -16px}.ZfdVuf .Y9aYob:focus:not(:hover)::before,.ZfdVuf .Y9aYob.u3bW4e::before{display:none}.ZfdVuf .Y9aYob:has(.GliO4d:focus-visible){--gm3-focus-ring-outward-display:block}.Y9aYob:empty,.XQ6hEf:empty{display:none}.uY2Qad{margin:0 0 24px}.ZfdVuf[data-expand-type="1"] .GliO4d{display:-webkit-box;display:-webkit-flex;display:flex}.ZfdVuf>.Y9aYob .xHr6Xe{-webkit-box-align:start;-webkit-align-items:flex-start;align-items:flex-start;padding-bottom:8px;padding-top:12px;position:relative;font-family:Google Sans,Roboto,Noto Sans Myanmar UI,Arial,sans-serif;font-weight:500;font-size:1rem;letter-spacing:0rem;line-height:1.5rem}.ZfdVuf:has(.XQ6hEf:empty)>.Y9aYob .xHr6Xe{padding-bottom:12px}.ySLakb.S7S4N .ySLakb .xHr6Xe{font-family:Google Sans,Roboto,Noto Sans Myanmar UI,Arial,sans-serif;font-weight:500;font-size:1rem;letter-spacing:0rem;line-height:1.5rem}.GliO4d{background:none;border:none;color:inherit;cursor:pointer;-webkit-box-flex:1;-webkit-flex-grow:1;flex-grow:1;font:inherit;margin:0;outline:0;padding:0;text-align:inherit}.GliO4d::-moz-focus-inner{border:0}.GliO4d .M0cpdd{color:var(--gm3-sys-color-on-surface,#1f1f1f);-webkit-box-flex:1;-webkit-flex-grow:1;flex-grow:1}.GliO4d .M0cpdd,.GliO4d .T5OKle{margin-top:4px}.h5Vxbc{-webkit-box-align:center;-webkit-align-items:center;align-items:center;background:var(--gm3-sys-color-secondary-container,#c2e7ff);border-radius:16px;color:var(--gm3-sys-color-on-secondary-container,#004a77);display:-webkit-box;display:-webkit-flex;display:flex;-webkit-flex-shrink:0;flex-shrink:0;height:32px;-webkit-box-pack:center;-webkit-justify-content:center;justify-content:center;margin-left:16px;width:28px}.h5Vxbc .kV7hid{-webkit-box-align:center;-webkit-align-items:center;align-items:center;display:-webkit-box;display:-webkit-flex;display:flex;height:20px;-webkit-box-pack:center;-webkit-justify-content:center;justify-content:center;-webkit-transition:-webkit-transform 0.2s cubic-bezier(0.4,0,0.2,1);transition:-webkit-transform 0.2s cubic-bezier(0.4,0,0.2,1);transition:transform 0.2s cubic-bezier(0.4,0,0.2,1);transition:transform 0.2s cubic-bezier(0.4,0,0.2,1),-webkit-transform 0.2s cubic-bezier(0.4,0,0.2,1);width:20px}.ZfdVuf.jVwmLb .h5Vxbc{background:var(--gm3-sys-color-surface-container,#f0f4f9);color:var(--gm3-sys-color-on-surface-variant,#444746)}.ZfdVuf.jVwmLb .kV7hid{-webkit-transform:rotate(-180deg);transform:rotate(-180deg)}.T5OKle{color:var(--gm3-sys-color-on-surface-variant,#444746);-webkit-flex-shrink:0;flex-shrink:0;height:24px;margin-right:16px;width:24px}.T5OKle .jLPeif{height:100%;width:100%}.i3HiPd .T5OKle{margin-top:0}.i3HiPd.sj692e .T5OKle{color:var(--gm3-sys-color-primary,#0b57d0)}.i3HiPd.Xq8bDe .T5OKle{color:var(--gm3-sys-color-error,#b3261e)}.i3HiPd.rNe0id .T5OKle{color:var(
    --wf-color-warning-icon,#f09d00
  )}.i3HiPd.YFdWic .T5OKle{height:48px;left:16px;position:absolute;top:16px;width:48px}.XQ6hEf{color:var(--gm3-sys-color-on-surface-variant,#444746);font-family:Google Sans,Roboto,Noto Sans Myanmar UI,Arial,sans-serif;font-weight:400;font-size:0.875rem;letter-spacing:0rem;line-height:1.25rem}.xe7Heb .XQ6hEf{margin-bottom:8px}.ZfdVuf .XQ6hEf{padding-bottom:16px}.Y9aYob:empty+.F4tG3e{margin-top:0}.F4tG3e{margin-bottom:16px;margin-top:4px}.Ci1RI>.F4tG3e{color:var(--gm3-sys-color-on-surface-variant,#444746);margin-bottom:0;margin-top:16px}.i3HiPd>.F4tG3e{margin-bottom:0;margin-top:0}.F4tG3e:only-child{margin-bottom:0;margin-top:0}.ZfdVuf>.F4tG3e{margin-top:0;overflow:hidden;-webkit-transition:0.2s cubic-bezier(0.4,0,0.2,1);transition:0.2s cubic-bezier(0.4,0,0.2,1)}.ySLakb.jVwmLb>.F4tG3e{margin-bottom:0;margin-top:0;max-height:0;opacity:0;visibility:hidden}.F4tG3e>[jsslot]>:first-child:not(.i3HiPd){margin-top:0;padding-top:0}.F4tG3e>[jsslot]>:last-child:not(.i3HiPd){margin-bottom:0;padding-bottom:0}.WXCwYb{display:none;margin-top:16px}.xe7Heb.jVwmLb .WXCwYb{display:block}.WXCwYb .hy0HVb{width:100%}.ySLakb.RDPZE{pointer-events:none}.ySLakb.RDPZE .xHr6Xe,.ySLakb.RDPZE .XQ6hEf,.ySLakb.RDPZE .F4tG3e,.ySLakb.RDPZE .T5OKle{color:var(--gm3-sys-color-on-surface,#1f1f1f);opacity:0.38}.jfyXNd .VfPpkd-IE5DDf{background-color:var(--gm3-sys-color-scrim,#000);opacity:0.32}.jfyXNd .VfPpkd-P5QLlc{background-color:var(--gm3-sys-color-surface-container-high,#e9eef6);border-radius:23px}.jfyXNd .VfPpkd-k2Wrsb{color:var(--gm3-sys-color-on-surface,#1f1f1f);font-family:Google Sans,Roboto,Noto Sans Myanmar UI,Arial,sans-serif;font-weight:400;font-size:1.5rem;letter-spacing:0rem;line-height:2rem}.jfyXNd .VfPpkd-cnG4Wd{color:var(--gm3-sys-color-on-surface-variant,#444746);padding-bottom:0;font-family:Google Sans,Roboto,Noto Sans Myanmar UI,Arial,sans-serif;font-weight:400;font-size:0.875rem;letter-spacing:0rem;line-height:1.25rem}.jfyXNd .VfPpkd-T0kwCb{padding:0 24px 16px 24px}.jfyXNd .F4tG3e{margin-left:0;margin-right:0;padding-left:0;padding-right:0}.jfyXNd .ksBjEc{color:var(--gm3-sys-color-primary,#0b57d0);font-size:0.875rem;height:40px;padding:0 16px}.jfyXNd .ksBjEc:hover:not(:disabled){color:var(--gm3-sys-color-primary,#0b57d0)}.jfyXNd .ksBjEc .VfPpkd-Jh9lGc::after,.jfyXNd .ksBjEc .VfPpkd-Jh9lGc::before{background-color:var(--gm3-sys-color-primary,#0b57d0)}.jfyXNd .ksBjEc:focus:not(:disabled){color:var(--gm3-sys-color-primary,#0b57d0)}.jfyXNd .ksBjEc .VfPpkd-J1Ukfc-LhBDec{border-color:var(--gm3-sys-color-primary,#0b57d0)}.jfyXNd .ksBjEc .VfPpkd-J1Ukfc-LhBDec::after{border-color:var(--gm3-sys-color-primary-container,#d3e3fd)}.jfyXNd .ksBjEc .VfPpkd-J1Ukfc-LhBDec::after,.jfyXNd .ksBjEc .VfPpkd-J1Ukfc-LhBDec,.jfyXNd .ksBjEc .VfPpkd-Jh9lGc{border-radius:23px}.jfyXNd.Zttm2{border-radius:0}.jfyXNd.Zttm2 .VfPpkd-P5QLlc{height:100vh;max-height:none;max-width:none;width:100vw}.jfyXNd.Zttm2 .yHy1rc{color:var(--gm3-sys-color-on-surface-variant,#444746);display:inline-block;padding:12px;text-align:center}.jfyXNd.Zttm2 .VfPpkd-zMU9ub .NMm5M{fill:var(--gm3-sys-color-primary,#0b57d0)}.jfyXNd.Zttm2 .VfPpkd-Bz112c-J1Ukfc-LhBDec{border-color:var(--gm3-sys-color-primary,#0b57d0);padding:2px}.jfyXNd.Zttm2 .VfPpkd-Bz112c-J1Ukfc-LhBDec,.jfyXNd.Zttm2 .VfPpkd-Bz112c-J1Ukfc-LhBDec::after{border-radius:50%}.jfyXNd.Zttm2 .yHy1rc:not(.VfPpkd-Bz112c-J1Ukfc-LhBDec)::before{display:none}.jfyXNd.Zttm2 .yHy1rc:not(.VfPpkd-Bz112c-J1Ukfc-LhBDec)::after{background:none;border:none;box-shadow:none}.jfyXNd.Zttm2 .yHy1rc .VfPpkd-Bz112c-Jh9lGc::before,.jfyXNd.Zttm2 .yHy1rc .VfPpkd-Bz112c-Jh9lGc::after{background-color:var(--gm3-sys-color-primary,#0b57d0)}.Zttm2 .qrsXKd{height:100%;width:100%}.Zttm2 .ToUTc{border:none;color-scheme:normal;display:block;height:100%;padding:0;width:100%}.qpGfHd{color:var(--gm3-sys-color-on-surface-variant,#444746);-webkit-box-flex:1;-webkit-flex-grow:1;flex-grow:1;padding-left:16px;font-family:Google Sans,Roboto,Noto Sans Myanmar UI,Arial,sans-serif;font-weight:400;font-size:0.875rem;letter-spacing:0rem;line-height:1.25rem}.XjS9D{display:-webkit-inline-box;display:-webkit-inline-flex;display:inline-flex}.XjS9D .VfPpkd-J1Ukfc-LhBDec{border-radius:22px}.XjS9D .VfPpkd-J1Ukfc-LhBDec::after{border-radius:24px}.XjS9D.eLNT1d{display:none}.XjS9D .TrZEUc .WpHeLc{position:absolute}.XjS9D.XjS9D .q6oraf .DMZ54e,.XjS9D.XjS9D .BqKGqe{font-family:"Google Sans",roboto,"Noto Sans Myanmar UI",arial,sans-serif;font-size:0.875rem;font-weight:500;font-weight:var(
    --c-afwt,500
  );letter-spacing:0rem;line-height:1.4285714286}.BqKGqe,.BqKGqe .VfPpkd-Jh9lGc{border-radius:20px}.XjS9D .VfPpkd-LgbsSe{height:40px}@media (orientation:landscape){.XjS9D .VfPpkd-LgbsSe{height:40px}}.Jskylb:not(:disabled){background:#0b57d0;color:#fff}.pIzcPc:not(:disabled),.eR0mzb:not(:disabled){color:#0b57d0;outline:#747775}.Jskylb.Jskylb.Jskylb:not(:disabled){background-color:var(--gm3-sys-color-primary,#0b57d0)}.Jskylb.Jskylb.Jskylb:not(:disabled){color:var(--gm3-sys-color-on-primary,#fff)}.Jskylb.Jskylb.Jskylb:not(:disabled):hover{color:var(--gm3-sys-color-on-primary,#fff)}.Jskylb.Jskylb.Jskylb:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.Jskylb.Jskylb.Jskylb:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:var(--gm3-sys-color-on-primary,#fff)}.Jskylb.Jskylb.Jskylb:not(:disabled):not(:disabled):active{color:var(--gm3-sys-color-on-primary,#fff)}.pIzcPc.pIzcPc.pIzcPc:not(:disabled){color:var(--gm3-sys-color-primary,#0b57d0)}.pIzcPc.pIzcPc.pIzcPc:not(:disabled):hover{color:var(--gm3-sys-color-primary,#0b57d0)}.pIzcPc.pIzcPc.pIzcPc:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.pIzcPc.pIzcPc.pIzcPc:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:var(--gm3-sys-color-primary,#0b57d0)}.pIzcPc.pIzcPc.pIzcPc .VfPpkd-Jh9lGc::before{background-color:var(--gm3-sys-color-primary,#0b57d0)}.pIzcPc.pIzcPc.pIzcPc .VfPpkd-Jh9lGc::after{background-color:var(--gm3-sys-color-primary,#0b57d0)}.pIzcPc.pIzcPc.pIzcPc:not(:disabled){border-color:var(--gm3-sys-color-outline,#747775)}.pIzcPc.pIzcPc.pIzcPc:not(:disabled):hover{border-color:var(--gm3-sys-color-outline,#747775)}.pIzcPc.pIzcPc.pIzcPc:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.pIzcPc.pIzcPc.pIzcPc:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{border-color:var(--gm3-sys-color-outline,#747775)}.pIzcPc.pIzcPc.pIzcPc:not(:disabled):active,.pIzcPc.pIzcPc.pIzcPc:not(:disabled):focus:active{border-color:var(--gm3-sys-color-outline,#747775)}.eR0mzb.eR0mzb.eR0mzb:not(:disabled){color:var(--gm3-sys-color-primary,#0b57d0)}.eR0mzb.eR0mzb.eR0mzb:not(:disabled):hover{color:var(--gm3-sys-color-primary,#0b57d0)}.eR0mzb.eR0mzb.eR0mzb:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.eR0mzb.eR0mzb.eR0mzb:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:var(--gm3-sys-color-primary,#0b57d0)}.eR0mzb.eR0mzb.eR0mzb .VfPpkd-Jh9lGc::before{background-color:var(--gm3-sys-color-primary,#0b57d0)}.eR0mzb.eR0mzb.eR0mzb .VfPpkd-Jh9lGc::after{background-color:var(--gm3-sys-color-primary,#0b57d0)}.AnSR9d.AnSR9d.AnSR9d:not(:disabled){background-color:var(--gm3-sys-color-secondary-container,#c2e7ff)}.AnSR9d.AnSR9d.AnSR9d:not(:disabled){color:var(--gm3-sys-color-on-secondary-container,#004a77)}.AnSR9d.AnSR9d.AnSR9d:not(:disabled):hover{color:var(--gm3-sys-color-on-secondary-container,#004a77)}.AnSR9d.AnSR9d.AnSR9d:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.AnSR9d.AnSR9d.AnSR9d:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:var(--gm3-sys-color-on-secondary-container,#004a77)}.AnSR9d.AnSR9d.AnSR9d:not(:disabled):not(:disabled):active{color:var(--gm3-sys-color-on-secondary-container,#004a77)}.eR0mzb.VfPpkd-LgbsSe{min-width:0}.eR0mzb.VfPpkd-LgbsSe{padding-left:16px;padding-right:16px}.H76ePc{margin:auto;max-width:380px;overflow:hidden;position:relative}.H76ePc .LbOduc{position:relative;text-align:center}.JQ5tlb{border-radius:50%;color:var(--gm3-sys-color-on-surface-variant,#444746);overflow:hidden}.pGzURd{line-height:1.4285714286}.lPxAeb{width:100%}.lPxAeb .JQ5tlb{-webkit-box-flex:0;-webkit-flex:none;flex:none;height:28px;margin-right:12px;width:28px}.lPxAeb .LbOduc,.VUfHYd .LbOduc{display:-webkit-box;display:-webkit-flex;display:flex;-webkit-box-align:center;-webkit-align-items:center;align-items:center}.lPxAeb .LbOduc{-webkit-box-pack:center;-webkit-justify-content:center;justify-content:center}.H76ePc .JQ5tlb{height:64px;margin:0 auto 8px;width:64px}.MnFlu{border-radius:50%;display:block}.lPxAeb .MnFlu,.lPxAeb .Qk3oof,.lPxAeb .uHLU0{max-height:100%;max-width:100%}.H76ePc .MnFlu,.H76ePc .Qk3oof,.H76ePc .uHLU0{height:64px;width:64px}.VUfHYd{height:24px}.VUfHYd .JQ5tlb{display:-webkit-box;display:-webkit-flex;display:flex;height:24px;margin-right:8px;min-width:24px}.VUfHYd .MnFlu,.VUfHYd .Qk3oof,.VUfHYd .uHLU0{color:var(--gm3-sys-color-on-surface-variant,#444746);height:24px;width:24px}.VUfHYd .DOLDDf{overflow:hidden}.lPxAeb .DOLDDf{-webkit-box-flex:1;-webkit-flex-grow:1;flex-grow:1}.lPxAeb .pGzURd{color:#1f1f1f;color:var(--gm3-sys-color-on-surface,#1f1f1f);font-family:"Google Sans",roboto,"Noto Sans Myanmar UI",arial,sans-serif;font-size:1rem;font-weight:500;letter-spacing:0rem;line-height:1.5}.H76ePc .pGzURd{color:#1f1f1f;color:var(--gm3-sys-color-on-surface,#1f1f1f);font-size:0.875rem}.yAlK0b,.VhdzSd,.H2oig{direction:ltr;font-size:0.875rem;line-height:1.4285714286;text-align:left;word-break:break-all}.yAlK0b{text-decoration:none}.lPxAeb .yAlK0b,.lPxAeb .VhdzSd,.lPxAeb .H2oig{font-size:0.875rem;font-weight:400;letter-spacing:0rem;line-height:1.4285714286}.H2oig{color:#444746;color:var(--gm3-sys-color-on-surface-variant,#444746)}.VUfHYd .yAlK0b{color:#1f1f1f;color:var(--gm3-sys-color-on-surface,#1f1f1f);font-family:"Google Sans",roboto,"Noto Sans Myanmar UI",arial,sans-serif;font-size:0.875rem;font-weight:500;letter-spacing:0rem;overflow:hidden;text-overflow:ellipsis;white-space:nowrap}.lPxAeb .VhdzSd{color:#444746;color:var(--gm3-sys-color-on-surface-variant,#444746)}.lPxAeb .yAlK0b{color:#444746;color:var(--gm3-sys-color-on-surface-variant,#444746)}.lPxAeb .yAlK0b[data-email$="@glimitedaccount.com"]{display:none}.H76ePc .yAlK0b{color:#444746;color:var(--gm3-sys-color-on-surface-variant,#444746)}.lrLKwc{color:#444746;color:var(--gm3-sys-color-on-surface-variant,#444746);font-size:0.875rem}.lPxAeb .lrLKwc{-webkit-align-self:flex-start;align-self:flex-start;-webkit-box-flex:0;-webkit-flex:none;flex:none;font-family:"Google Sans",roboto,"Noto Sans Myanmar UI",arial,sans-serif;font-size:0.75rem;font-weight:400;letter-spacing:0.00625rem;line-height:1.3333333333}.Ahygpe{-webkit-box-align:center;-webkit-align-items:center;align-items:center;background:#fff;background:var(--gm3-sys-color-surface-container-lowest,#fff);border:1px solid var(--gm3-sys-color-outline,#747775);color:var(--gm3-sys-color-on-surface,#1f1f1f);cursor:pointer;display:-webkit-inline-box;display:-webkit-inline-flex;display:inline-flex;font-size:0.875rem;font-weight:500;letter-spacing:.25px;max-width:100%;position:relative}.Ahygpe::after{border:1px solid transparent;content:"";position:absolute;inset:-1px}.Ahygpe:focus-visible::after{border:2px solid;border-color:#0b57d0;border-color:var(--gm3-sys-color-primary,#0b57d0);box-shadow:0 0 0 2px #d3e3fd;box-shadow:0 0 0 2px var(--gm3-sys-color-primary-container,#d3e3fd);border-radius:26px;content:"";position:absolute;pointer-events:none;inset:-5px}.Zjyti{color:#0b57d0;color:var(--gm3-sys-color-primary,#0b57d0);font-size:0.75rem}.m8wwGd{border-radius:16px;padding:0 15px 0 15px}.m8wwGd{position:relative}.m8wwGd::before{background:#1f1f1f;background:var(--gm3-sys-color-on-surface,#1f1f1f);content:"";opacity:0;position:absolute;pointer-events:none}.m8wwGd:hover::before{opacity:0.08}.m8wwGd:focus::before,.m8wwGd.u3bW4e::before{opacity:0.1}.m8wwGd:active::before,.m8wwGd.qs41qe::before{opacity:0.1}.m8wwGd::before{border-radius:16px;width:100%;height:100%}.m8wwGd:focus,.m8wwGd.u3bW4e{outline:none;border-color:#747775;border-color:var(--gm3-sys-color-outline,#747775)}.m8wwGd:active,.m8wwGd.qs41qe{color:#1f1f1f;color:var(--gm3-sys-color-on-surface,#1f1f1f);border-color:#1f1f1f;border-color:var(--gm3-sys-color-on-surface,#1f1f1f)}.m8wwGd.Zjyti{border-radius:12px;padding:0 10px 0 10px}.m8wwGd.EPPJc{padding-right:8px}.m8wwGd.cd29Sd{padding-left:3px}.m8wwGd.Zjyti.EPPJc{padding-right:8px}.m8wwGd.Zjyti.cd29Sd{padding-left:2px}.m8wwGd::after{border-radius:16px}.m8wwGd.Zjyti::after{border-radius:12px}.HOE91e{border-radius:12px;height:24px;margin-right:8px}.HOE91e .MnFlu,.HOE91e .Qk3oof,.HOE91e .uHLU0{border-radius:50%;color:var(--gm3-sys-color-on-surface-variant,#444746);display:block;height:24px;width:24px}.IxcUte{direction:ltr;text-align:left;overflow:hidden;text-overflow:ellipsis;white-space:nowrap}.m8wwGd .IxcUte{line-height:30px}.m8wwGd.xNLKcb .IxcUte{font-family:"Google Sans",roboto,"Noto Sans Myanmar UI",arial,sans-serif;font-size:0.875rem;font-weight:500;letter-spacing:0rem;text-decoration:none}.m8wwGd.Zjyti .IxcUte{line-height:22px}.JCl8ie{color:var(--gm3-sys-color-on-surface,#1f1f1f);-webkit-flex-shrink:0;flex-shrink:0;height:20px;margin-left:5px;width:20px;-webkit-transition:-webkit-transform 0.2s cubic-bezier(0.4,0,0.2,1);transition:-webkit-transform 0.2s cubic-bezier(0.4,0,0.2,1);transition:transform 0.2s cubic-bezier(0.4,0,0.2,1);transition:transform 0.2s cubic-bezier(0.4,0,0.2,1),-webkit-transform 0.2s cubic-bezier(0.4,0,0.2,1)}.Ahygpe.sMVRZe .JCl8ie{-webkit-transform:rotate(180deg);transform:rotate(180deg)}.Zjyti .JCl8ie{height:16px;width:16px}.u4TTuf{display:block;height:100%;width:100%}.rFrNMe{-webkit-user-select:none;-webkit-user-select:none;-webkit-tap-highlight-color:transparent;display:inline-block;outline:none;padding-bottom:8px;width:200px}.aCsJod{height:40px;position:relative;vertical-align:top}.aXBtI{display:-webkit-box;display:-webkit-flex;display:-webkit-box;display:-webkit-flex;display:flex;position:relative;top:14px}.Xb9hP{display:-webkit-box;display:-webkit-flex;display:-webkit-box;display:-webkit-flex;display:flex;-webkit-box-flex:1;-webkit-flex-grow:1;-webkit-box-flex:1;box-flex:1;-webkit-flex-grow:1;flex-grow:1;-webkit-flex-shrink:1;-webkit-flex-shrink:1;flex-shrink:1;min-width:0%;position:relative}.A37UZe{-webkit-box-sizing:border-box;box-sizing:border-box;height:24px;line-height:24px;position:relative}.qgcB3c:not(:empty){padding-right:12px}.sxyYjd:not(:empty){padding-left:12px}.whsOnd{-webkit-box-flex:1;-webkit-flex-grow:1;-webkit-box-flex:1;box-flex:1;-webkit-flex-grow:1;flex-grow:1;-webkit-flex-shrink:1;-webkit-flex-shrink:1;flex-shrink:1;background-color:transparent;border:none;display:block;font:400 16px Roboto,RobotoDraft,Helvetica,Arial,sans-serif;height:24px;line-height:24px;margin:0;min-width:0%;outline:none;padding:0;z-index:0}.rFrNMe.dm7YTc .whsOnd{color:#fff}.whsOnd:invalid,.whsOnd:-moz-submit-invalid,.whsOnd:-moz-ui-invalid{-webkit-box-shadow:none;box-shadow:none}.I0VJ4d>.whsOnd::-ms-clear,.I0VJ4d>.whsOnd::-ms-reveal{display:none}.i9lrp{background-color:rgba(0,0,0,.12);bottom:-2px;height:1px;left:0;margin:0;padding:0;position:absolute;width:100%}.i9lrp::before{content:"";position:absolute;top:0;bottom:-2px;left:0;right:0;border-bottom:1px solid rgba(0,0,0,0);pointer-events:none}.rFrNMe.dm7YTc .i9lrp{background-color:rgba(255,255,255,.7)}.OabDMe{-webkit-transform:scaleX(0);-webkit-transform:scaleX(0);transform:scaleX(0);background-color:#4285f4;bottom:-2px;height:2px;left:0;margin:0;padding:0;position:absolute;width:100%}.rFrNMe.dm7YTc .OabDMe{background-color:#a1c2fa}.rFrNMe.k0tWj .i9lrp,.rFrNMe.k0tWj .OabDMe{background-color:#d50000;height:2px}.rFrNMe.k0tWj.dm7YTc .i9lrp,.rFrNMe.k0tWj.dm7YTc .OabDMe{background-color:#e06055}.whsOnd[disabled]{color:rgba(0,0,0,.38)}.rFrNMe.dm7YTc .whsOnd[disabled]{color:rgba(255,255,255,.5)}.whsOnd[disabled]~.i9lrp{background:none;border-bottom:1px dotted rgba(0,0,0,.38)}.OabDMe.Y2Zypf{-webkit-animation:quantumWizPaperInputRemoveUnderline .3s cubic-bezier(0.4,0,0.2,1);-webkit-animation:quantumWizPaperInputRemoveUnderline .3s cubic-bezier(0.4,0,0.2,1);animation:quantumWizPaperInputRemoveUnderline .3s cubic-bezier(0.4,0,0.2,1)}.rFrNMe.u3bW4e .OabDMe{-webkit-animation:quantumWizPaperInputAddUnderline .3s cubic-bezier(0.4,0,0.2,1);-webkit-animation:quantumWizPaperInputAddUnderline .3s cubic-bezier(0.4,0,0.2,1);animation:quantumWizPaperInputAddUnderline .3s cubic-bezier(0.4,0,0.2,1);-webkit-transform:scaleX(1);-webkit-transform:scaleX(1);transform:scaleX(1)}.rFrNMe.sdJrJc>.aCsJod{padding-top:24px}.AxOyFc{-webkit-transform-origin:bottom left;-webkit-transform-origin:bottom left;transform-origin:bottom left;-webkit-transition:all .3s cubic-bezier(0.4,0,0.2,1);-webkit-transition:all .3s cubic-bezier(0.4,0,0.2,1);transition:all .3s cubic-bezier(0.4,0,0.2,1);-webkit-transition-property:color,bottom,-webkit-transform;-webkit-transition-property:color,bottom,-webkit-transform;transition-property:color,bottom,-webkit-transform;-webkit-transition-property:color,bottom,transform;transition-property:color,bottom,transform;-webkit-transition-property:color,bottom,transform,-webkit-transform;transition-property:color,bottom,transform,-webkit-transform;color:rgba(0,0,0,.38);font:400 16px Roboto,RobotoDraft,Helvetica,Arial,sans-serif;font-size:16px;pointer-events:none;position:absolute;bottom:3px;left:0;width:100%}.whsOnd:not([disabled]):focus~.AxOyFc,.whsOnd[badinput=true]~.AxOyFc,.rFrNMe.CDELXb .AxOyFc,.rFrNMe.dLgj8b .AxOyFc{-webkit-transform:scale(0.75) translateY(-39px);-webkit-transform:scale(0.75) translateY(-39px);transform:scale(0.75) translateY(-39px)}.whsOnd:not([disabled]):focus~.AxOyFc{color:#3367d6}.rFrNMe.dm7YTc .whsOnd:not([disabled]):focus~.AxOyFc{color:#a1c2fa}.rFrNMe.k0tWj .whsOnd:not([disabled]):focus~.AxOyFc{color:#d50000}.ndJi5d{color:rgba(0,0,0,.38);font:400 16px Roboto,RobotoDraft,Helvetica,Arial,sans-serif;max-width:100%;overflow:hidden;pointer-events:none;position:absolute;text-overflow:ellipsis;top:2px;left:0;white-space:nowrap}.rFrNMe.CDELXb .ndJi5d{display:none}.K0Y8Se{-webkit-tap-highlight-color:transparent;font:400 12px Roboto,RobotoDraft,Helvetica,Arial,sans-serif;height:16px;margin-left:auto;padding-left:16px;padding-top:8px;pointer-events:none;opacity:.3;white-space:nowrap}.rFrNMe.dm7YTc .AxOyFc,.rFrNMe.dm7YTc .K0Y8Se,.rFrNMe.dm7YTc .ndJi5d{color:rgba(255,255,255,.7)}.rFrNMe.Tyc9J{padding-bottom:4px}.dEOOab,.ovnfwe:not(:empty){-webkit-tap-highlight-color:transparent;-webkit-box-flex:1;-webkit-flex:1 1 auto;-webkit-box-flex:1 1 auto;-webkit-flex:1 1 auto;flex:1 1 auto;font:400 12px Roboto,RobotoDraft,Helvetica,Arial,sans-serif;min-height:16px;padding-top:8px}.LXRPh{display:-webkit-box;display:-webkit-flex;display:-webkit-box;display:-webkit-flex;display:flex}.ovnfwe{pointer-events:none}.dEOOab{color:#d50000}.rFrNMe.dm7YTc .dEOOab,.rFrNMe.dm7YTc.k0tWj .whsOnd:not([disabled]):focus~.AxOyFc{color:#e06055}.ovnfwe{opacity:.3}.rFrNMe.dm7YTc .ovnfwe{color:rgba(255,255,255,.7);opacity:1}.rFrNMe.k0tWj .ovnfwe,.rFrNMe:not(.k0tWj) .ovnfwe:not(:empty)+.dEOOab{display:none}@-webkit-keyframes quantumWizPaperInputRemoveUnderline{0%{-webkit-transform:scaleX(1);-webkit-transform:scaleX(1);transform:scaleX(1);opacity:1}to{-webkit-transform:scaleX(1);-webkit-transform:scaleX(1);transform:scaleX(1);opacity:0}}@keyframes quantumWizPaperInputRemoveUnderline{0%{-webkit-transform:scaleX(1);-webkit-transform:scaleX(1);transform:scaleX(1);opacity:1}to{-webkit-transform:scaleX(1);-webkit-transform:scaleX(1);transform:scaleX(1);opacity:0}}@-webkit-keyframes quantumWizPaperInputAddUnderline{0%{-webkit-transform:scaleX(0);-webkit-transform:scaleX(0);transform:scaleX(0)}to{-webkit-transform:scaleX(1);-webkit-transform:scaleX(1);transform:scaleX(1)}}@keyframes quantumWizPaperInputAddUnderline{0%{-webkit-transform:scaleX(0);-webkit-transform:scaleX(0);transform:scaleX(0)}to{-webkit-transform:scaleX(1);-webkit-transform:scaleX(1);transform:scaleX(1)}}@media (min-width:600px){.njnYzb.DbQnIe .YqLCIe{display:-webkit-box;display:-webkit-flex;display:flex;-webkit-box-pack:justify;-webkit-justify-content:space-between;justify-content:space-between}}.njnYzb:first-child .H2p7Gf:first-child .i79UJc{padding-top:8px}@media (min-width:600px){.njnYzb.DbQnIe:first-child .H2p7Gf .i79UJc{padding-top:8px}.njnYzb.DbQnIe .H2p7Gf{-webkit-box-flex:1;-webkit-flex-grow:1;flex-grow:1;margin-right:8px;width:0}.njnYzb.DbQnIe .H2p7Gf:last-child{margin-right:0}}.i79UJc.i79UJc{box-sizing:content-box}.i79UJc{padding-bottom:0;padding-top:24px;width:100%}.i79UJc .oJeWuf.oJeWuf{height:56px;padding-top:0}.i79UJc.OcVpRe .oJeWuf.oJeWuf{height:36px}.i79UJc .Wic03c{-webkit-box-align:center;-webkit-align-items:center;align-items:center;position:static}.i79UJc .snByac{background-color:transparent;bottom:18px;box-sizing:border-box;color:var(--gm3-sys-color-on-surface-variant,#444746);font-size:16px;font-weight:400;left:8px;max-width:calc(100% - 16px);overflow:hidden;padding:0 8px;text-overflow:ellipsis;-webkit-transition:opacity .15s cubic-bezier(.4,0,.2,1),background-color .15s cubic-bezier(.4,0,.2,1),-webkit-transform .15s cubic-bezier(.4,0,.2,1);transition:opacity .15s cubic-bezier(.4,0,.2,1),background-color .15s cubic-bezier(.4,0,.2,1),-webkit-transform .15s cubic-bezier(.4,0,.2,1);transition:transform .15s cubic-bezier(.4,0,.2,1),opacity .15s cubic-bezier(.4,0,.2,1),background-color .15s cubic-bezier(.4,0,.2,1);transition:transform .15s cubic-bezier(.4,0,.2,1),opacity .15s cubic-bezier(.4,0,.2,1),background-color .15s cubic-bezier(.4,0,.2,1),-webkit-transform .15s cubic-bezier(.4,0,.2,1);white-space:nowrap;width:auto;z-index:1}.i79UJc.OcVpRe .snByac{bottom:10px;color:var(--gm3-sys-color-on-surface-variant,#444746);font-size:14px;left:4px;line-height:16px;padding:0 6px}.i79UJc.u3bW4e .snByac.snByac,.i79UJc.CDELXb .snByac.snByac{background-color:#fff;background-color:var(--gm3-sys-color-surface-container-lowest,#fff);-webkit-transform:scale(.75) translatey(-41px);transform:scale(.75) translatey(-41px)}.i79UJc.OcVpRe.u3bW4e .snByac,.i79UJc.OcVpRe.CDELXb .snByac{-webkit-transform:scale(.75) translatey(-165%);transform:scale(.75) translatey(-165%)}.i79UJc .zHQkBf:not([disabled]):focus~.snByac{color:#0b57d0;color:var(--gm3-sys-color-primary,#0b57d0)}.i79UJc.IYewr.u3bW4e .zHQkBf:not([disabled])~.snByac,.i79UJc.IYewr.CDELXb .zHQkBf:not([disabled])~.snByac{color:#b3261e;color:var(--gm3-sys-color-error,#b3261e)}.i79UJc .zHQkBf{border-radius:4px;color:#1f1f1f;color:var(--gm3-sys-color-on-surface,#1f1f1f);font-family:"Google Sans",roboto,"Noto Sans Myanmar UI",arial,sans-serif;font-size:16px;height:28px;margin:2px;padding:12px 14px;text-align:left;z-index:1}.i79UJc.OcVpRe .zHQkBf{font-size:14px;height:20px;padding:6px 8px}.i79UJc.YKooDc .zHQkBf,.i79UJc.YKooDc .MQL3Ob{direction:ltr;text-align:left}.i79UJc .iHd5yb{padding-left:14px}.i79UJc.OcVpRe .iHd5yb{padding-left:8px}.i79UJc .MQL3Ob{padding-right:14px;z-index:1}.i79UJc.OcVpRe .MQL3Ob{padding-right:8px}.i79UJc .mIZh1c,.i79UJc .cXrdqd{border-radius:4px;bottom:0;box-sizing:border-box}.i79UJc .mIZh1c,.i79UJc .cXrdqd,.i79UJc.IYewr .mIZh1c,.i79UJc.IYewr .cXrdqd{background-color:transparent;bottom:0;height:auto;top:0}.i79UJc .mIZh1c{border:1px solid;border-color:#747775;border-color:var(--gm3-sys-color-outline,#747775);padding:1px}.i79UJc .cXrdqd{border:1px solid;border-color:#0b57d0;border-color:var(--gm3-sys-color-primary,#0b57d0);opacity:0;-webkit-transform:none;transform:none;-webkit-transition:opacity .15s cubic-bezier(.4,0,.2,1);transition:opacity .15s cubic-bezier(.4,0,.2,1)}.i79UJc.u3bW4e .cXrdqd{border-width:2px}.i79UJc.u3bW4e .cXrdqd,.i79UJc.IYewr .cXrdqd{-webkit-animation:none;animation:none;opacity:1}.i79UJc.IYewr .cXrdqd{border-color:#b3261e;border-color:var(--gm3-sys-color-error,#b3261e)}.i79UJc .ndJi5d,.i79UJc .ovnfwe{pointer-events:auto}.i79UJc .RxsGPe,.i79UJc .Is7Fhb{display:none}.Ly8vae{color:#444746;color:var(--gm3-sys-color-on-surface-variant,#444746);display:-webkit-box;display:-webkit-flex;display:flex;font-family:"Google Sans",roboto,"Noto Sans Myanmar UI",arial,sans-serif;font-size:0.75rem;font-weight:400;letter-spacing:0.00625rem;line-height:1.3333333333}.Ly8vae:empty,.NdBX9e:empty{display:none}.njnYzb.Jj6Lae .Ly8vae{color:#b3261e;color:var(--gm3-sys-color-error,#b3261e)}.jEOsLc{display:none;margin-right:8px}.JPqhye{height:16px;width:16px}.njnYzb.Jj6Lae .jEOsLc{display:block}.njnYzb .Ly8vae{color:#444746;color:var(--gm3-sys-color-on-surface-variant,#444746);margin-top:4px}.njnYzb .YQOsOe{margin-left:16px}.njnYzb.OcVpRe .YQOsOe{margin-left:10px}.Ekjuhf{color:#444746;color:var(--gm3-sys-color-on-surface-variant,#444746);-webkit-box-align:start;-webkit-align-items:flex-start;align-items:flex-start;display:-webkit-box;display:-webkit-flex;display:flex;font-family:"Google Sans",roboto,"Noto Sans Myanmar UI",arial,sans-serif;font-size:0.75rem;font-weight:400;letter-spacing:0.00625rem;line-height:1.3333333333;margin-top:2px}.Ekjuhf.Jj6Lae{color:#b3261e;color:var(--gm3-sys-color-error,#b3261e)}.AfGCob{margin-right:8px;margin-top:calc((1px*var(--boq-accounts-wireframe-themes-materialnext-common-abstractinput-help-line-height-unitless-px) - 16px)/2)}.xTjuxe{display:block;height:16px;width:16px}.edhGSc{-webkit-user-select:none;-webkit-user-select:none;-webkit-tap-highlight-color:transparent;display:inline-block;outline:none;padding-bottom:8px}.RpC4Ne{min-height:1.5em;position:relative;vertical-align:top}.Pc9Gce{display:-webkit-box;display:-webkit-flex;display:-webkit-box;display:-webkit-flex;display:flex;position:relative;padding-top:14px}.KHxj8b{-webkit-box-flex:1;-webkit-flex-grow:1;-webkit-box-flex:1;box-flex:1;-webkit-flex-grow:1;flex-grow:1;-webkit-flex-shrink:1;-webkit-flex-shrink:1;flex-shrink:1;background-color:transparent;border:none;display:block;font:400 16px Roboto,RobotoDraft,Helvetica,Arial,sans-serif;height:24px;min-height:24px;line-height:24px;margin:0;outline:none;padding:0;resize:none;white-space:pre-wrap;word-wrap:break-word;z-index:0;overflow-y:visible;overflow-x:hidden}.KHxj8b.VhWN2c{text-align:center}.edhGSc.dm7YTc .KHxj8b{color:rgba(255,255,255,.87)}.edhGSc.u3bW4e.dm7YTc .KHxj8b{color:#fff}.z0oSpf{background-color:rgba(0,0,0,.12);height:1px;left:0;margin:0;padding:0;position:absolute;width:100%}.edhGSc.dm7YTc>.RpC4Ne>.z0oSpf{background-color:rgba(255,255,255,.12)}.Bfurwb{-webkit-transform:scaleX(0);-webkit-transform:scaleX(0);transform:scaleX(0);background-color:#4285f4;height:2px;left:0;margin:0;padding:0;position:absolute;width:100%}.edhGSc.k0tWj>.RpC4Ne>.z0oSpf,.edhGSc.k0tWj>.RpC4Ne>.Bfurwb{background-color:#d50000;height:2px}.edhGSc.k0tWj.dm7YTc>.RpC4Ne>.z0oSpf,.edhGSc.k0tWj.dm7YTc>.RpC4Ne>.Bfurwb{background-color:#ff6e6e}.edhGSc.RDPZE .KHxj8b{color:rgba(0,0,0,.38)}.edhGSc.RDPZE>.RpC4Ne>.z0oSpf{background:none;border-bottom:1px dotted rgba(0,0,0,.38)}.Bfurwb.Y2Zypf{-webkit-animation:quantumWizPaperInputRemoveUnderline .3s cubic-bezier(0.4,0,0.2,1);-webkit-animation:quantumWizPaperInputRemoveUnderline .3s cubic-bezier(0.4,0,0.2,1);animation:quantumWizPaperInputRemoveUnderline .3s cubic-bezier(0.4,0,0.2,1)}.edhGSc.u3bW4e>.RpC4Ne>.Bfurwb{-webkit-animation:quantumWizPaperInputAddUnderline .3s cubic-bezier(0.4,0,0.2,1);-webkit-animation:quantumWizPaperInputAddUnderline .3s cubic-bezier(0.4,0,0.2,1);animation:quantumWizPaperInputAddUnderline .3s cubic-bezier(0.4,0,0.2,1);-webkit-transform:scaleX(1);-webkit-transform:scaleX(1);transform:scaleX(1)}.edhGSc.FPYHkb>.RpC4Ne{padding-top:24px}.fqp6hd{-webkit-transform-origin:top left;-webkit-transform-origin:top left;transform-origin:top left;-webkit-transform:translate(0,-22px);-webkit-transform:translate(0,-22px);transform:translate(0,-22px);-webkit-transition:all .3s cubic-bezier(0.4,0,0.2,1);-webkit-transition:all .3s cubic-bezier(0.4,0,0.2,1);transition:all .3s cubic-bezier(0.4,0,0.2,1);-webkit-transition-property:color,top,-webkit-transform;-webkit-transition-property:color,top,-webkit-transform;transition-property:color,top,-webkit-transform;-webkit-transition-property:color,top,transform;transition-property:color,top,transform;-webkit-transition-property:color,top,transform,-webkit-transform;transition-property:color,top,transform,-webkit-transform;color:rgba(0,0,0,.38);font:400 16px Roboto,RobotoDraft,Helvetica,Arial,sans-serif;font-size:16px;pointer-events:none;position:absolute;top:100%;width:100%}.edhGSc.u3bW4e>.RpC4Ne>.fqp6hd,.edhGSc.CDELXb>.RpC4Ne>.fqp6hd,.edhGSc.LydCob .fqp6hd{-webkit-transform:scale(0.75);-webkit-transform:scale(0.75);transform:scale(0.75);top:16px}.edhGSc.dm7YTc>.RpC4Ne>.fqp6hd{color:rgba(255,255,255,.38)}.edhGSc.u3bW4e>.RpC4Ne>.fqp6hd,.edhGSc.u3bW4e.dm7YTc>.RpC4Ne>.fqp6hd{color:#4285f4}.F1pOBe{color:rgba(0,0,0,.38);font:400 16px Roboto,RobotoDraft,Helvetica,Arial,sans-serif;max-width:100%;overflow:hidden;pointer-events:none;position:absolute;bottom:3px;text-overflow:ellipsis;white-space:nowrap}.edhGSc.dm7YTc .F1pOBe{color:rgba(255,255,255,.38)}.edhGSc.CDELXb>.RpC4Ne>.F1pOBe{display:none}.S1BUyf{-webkit-tap-highlight-color:transparent;font:400 12px Roboto,RobotoDraft,Helvetica,Arial,sans-serif;height:16px;margin-left:auto;padding-left:16px;padding-top:8px;pointer-events:none;text-align:right;color:rgba(0,0,0,.38);white-space:nowrap}.edhGSc.dm7YTc>.S1BUyf{color:rgba(255,255,255,.38)}.edhGSc.wrxyb{padding-bottom:4px}.v6odTb,.YElZX:not(:empty){-webkit-tap-highlight-color:transparent;-webkit-box-flex:1;-webkit-flex:1 1 auto;-webkit-box-flex:1 1 auto;-webkit-flex:1 1 auto;flex:1 1 auto;font:400 12px Roboto,RobotoDraft,Helvetica,Arial,sans-serif;min-height:16px;padding-top:8px}.edhGSc.wrxyb .jE8NUc{display:-webkit-box;display:-webkit-flex;display:-webkit-box;display:-webkit-flex;display:flex}.YElZX{pointer-events:none}.v6odTb{color:#d50000}.edhGSc.dm7YTc .v6odTb{color:#ff6e6e}.YElZX{opacity:.3}.edhGSc.k0tWj .YElZX,.edhGSc:not(.k0tWj) .YElZX:not(:empty)+.v6odTb{display:none}@-webkit-keyframes quantumWizPaperInputRemoveUnderline{0%{-webkit-transform:scaleX(1);-webkit-transform:scaleX(1);transform:scaleX(1);opacity:1}to{-webkit-transform:scaleX(1);-webkit-transform:scaleX(1);transform:scaleX(1);opacity:0}}@keyframes quantumWizPaperInputRemoveUnderline{0%{-webkit-transform:scaleX(1);-webkit-transform:scaleX(1);transform:scaleX(1);opacity:1}to{-webkit-transform:scaleX(1);-webkit-transform:scaleX(1);transform:scaleX(1);opacity:0}}@-webkit-keyframes quantumWizPaperInputAddUnderline{0%{-webkit-transform:scaleX(0);-webkit-transform:scaleX(0);transform:scaleX(0)}to{-webkit-transform:scaleX(1);-webkit-transform:scaleX(1);transform:scaleX(1)}}@keyframes quantumWizPaperInputAddUnderline{0%{-webkit-transform:scaleX(0);-webkit-transform:scaleX(0);transform:scaleX(0)}to{-webkit-transform:scaleX(1);-webkit-transform:scaleX(1);transform:scaleX(1)}}.X3mtXb{box-sizing:content-box}.FAiUob,.X3mtXb{display:block;padding:16px 0 0;width:100%}.AFTWye.OcVpRe .X3mtXb,.AFTWye.OcVpRe .FAiUob{padding:24px 0 0;padding-bottom:0}:first-child>.X3mtXb,:first-child>.FAiUob,:first-child.OcVpRe>.X3mtXb,:first-child.OcVpRe>.FAiUob{padding:8px 0 0}.AFTWye .X3mtXb .oJeWuf{height:56px;padding-top:0}.AFTWye.OcVpRe .X3mtXb .oJeWuf{height:36px}.X3mtXb .Wic03c{-webkit-box-align:center;-webkit-align-items:center;align-items:center;position:static;top:0}.X3mtXb .snByac{background:#fff;background:var(--gm3-sys-color-surface-container-lowest,#fff);color:#444746;color:var(--gm3-sys-color-on-surface-variant,#444746);bottom:17px;box-sizing:border-box;font-size:16px;font-weight:400;left:8px;max-width:calc(100% - 16px);overflow:hidden;padding:0 8px;text-overflow:ellipsis;-webkit-transition:opacity .15s cubic-bezier(.4,0,.2,1),-webkit-transform .15s cubic-bezier(.4,0,.2,1);transition:opacity .15s cubic-bezier(.4,0,.2,1),-webkit-transform .15s cubic-bezier(.4,0,.2,1);transition:transform .15s cubic-bezier(.4,0,.2,1),opacity .15s cubic-bezier(.4,0,.2,1);transition:transform .15s cubic-bezier(.4,0,.2,1),opacity .15s cubic-bezier(.4,0,.2,1),-webkit-transform .15s cubic-bezier(.4,0,.2,1);white-space:nowrap;width:auto;z-index:1}.X3mtXb.IYewr.u3bW4e .zHQkBf:not([disabled])~.snByac{color:#b3261e;color:var(--gm3-sys-color-error,#b3261e)}.AFTWye.OcVpRe .X3mtXb .snByac{color:#444746;color:var(--gm3-sys-color-on-surface-variant,#444746);bottom:9px;font-size:14px;left:4px;line-height:16px;padding:0 6px}.AFTWye.OcVpRe .u3bW4e .snByac,.AFTWye.OcVpRe .CDELXb .snByac{-webkit-transform:scale(.75) translateY(-155%);transform:scale(.75) translateY(-155%)}.X3mtXb .ndJi5d{top:inherit}.X3mtXb .ndJi5d,.X3mtXb .ovnfwe{pointer-events:auto}.X3mtXb .Is7Fhb,.X3mtXb .RxsGPe{font-family:"Google Sans",roboto,"Noto Sans Myanmar UI",arial,sans-serif;font-size:0.75rem;font-weight:400;letter-spacing:0.00625rem;line-height:1.3333333333;opacity:1;padding-top:4px}.AFTWye .Is7Fhb{color:var(--gm3-sys-color-on-surface-variant,#444746);margin-left:16px}.AFTWye.OcVpRe .Is7Fhb{margin-left:10px}.X3mtXb .RxsGPe{color:#b3261e;color:var(--gm3-sys-color-error,#b3261e)}.X3mtXb .Is7Fhb:empty,.X3mtXb .RxsGPe:empty{display:none}.X3mtXb .zHQkBf{border-radius:4px;color:#1f1f1f;color:var(--gm3-sys-color-on-surface,#1f1f1f);font-family:"Google Sans",roboto,"Noto Sans Myanmar UI",arial,sans-serif;font-size:16px;height:28px;margin:1px 1px 0 1px;padding:13px 15px;text-align:left;width:100%;z-index:1}.X3mtXb.u3bW4e .zHQkBf,.X3mtXb.IYewr .zHQkBf{margin:2px 2px 0 2px;padding:12px 14px}.AFTWye.OcVpRe .X3mtXb .zHQkBf{font-size:14px;height:20px;padding:7px 9px}.AFTWye.OcVpRe .u3bW4e .zHQkBf,.AFTWye.OcVpRe .IYewr .zHQkBf{height:20px;padding:6px 8px}.UOsO2 .Wic03c,.UOsO2 .zHQkBf,.UOsO2 .iHd5yb,.UOsO2 .MQL3Ob{direction:ltr;text-align:left}.UOsO2 .Wic03c .snByac{direction:ltr}.X3mtXb .iHd5yb{padding-left:15px}.X3mtXb.u3bW4e .iHd5yb{padding-left:14px}.X3mtXb .MQL3Ob{padding-right:15px;z-index:1}.X3mtXb.u3bW4e .MQL3Ob{padding-right:15px}.AFTWye.OcVpRe .X3mtXb .iHd5yb{padding-left:9px}.AFTWye.OcVpRe .X3mtXb.u3bW4e .iHd5yb{padding-left:8px}.AFTWye.OcVpRe .X3mtXb .MQL3Ob,.AFTWye.OcVpRe .X3mtXb.u3bW4e .MQL3Ob{padding-right:9px}.X3mtXb .AxOyFc{font-family:"Google Sans",roboto,"Noto Sans Myanmar UI",arial,sans-serif}.X3mtXb .whsOnd:not([disabled]):focus~.AxOyFc{color:#0b57d0;color:var(--gm3-sys-color-primary,#0b57d0)}.X3mtXb .mIZh1c{border:1px solid;border-color:#747775;border-color:var(--gm3-sys-color-outline,#747775);border-radius:4px;bottom:0;box-sizing:border-box}.X3mtXb .cXrdqd{border-radius:4px;bottom:0;opacity:0;-webkit-transform:none;transform:none;-webkit-transition:opacity .15s cubic-bezier(.4,0,.2,1);transition:opacity .15s cubic-bezier(.4,0,.2,1);width:calc(100% - 4px)}.X3mtXb .mIZh1c,.X3mtXb .cXrdqd,.X3mtXb.IYewr .mIZh1c,.X3mtXb.IYewr .cXrdqd{background-color:transparent}.X3mtXb .mIZh1c,.X3mtXb.k0tWj .mIZh1c{height:100%}.X3mtXb.IYewr .cXrdqd{height:calc(100% - 2px);width:calc(100% - 2px)}.X3mtXb .cXrdqd,.X3mtXb.IYewr.u3bW4e .cXrdqd{height:calc(100% - 4px);width:calc(100% - 4px)}.X3mtXb.u3bW4e .cXrdqd,.X3mtXb.IYewr .cXrdqd{-webkit-animation:none;animation:none;opacity:1}.X3mtXb.u3bW4e .cXrdqd{border:2px solid;border-color:#0b57d0;border-color:var(--gm3-sys-color-primary,#0b57d0)}.X3mtXb.IYewr.u3bW4e .cXrdqd{border-width:2px}.X3mtXb.IYewr .cXrdqd{border:1px solid;border-color:#b3261e;border-color:var(--gm3-sys-color-error,#b3261e)}.X3mtXb.IYewr.CDELXb .snByac{color:#b3261e;color:var(--gm3-sys-color-error,#b3261e)}.X3mtXb .zHQkBf[disabled]{color:#1f1f1f;color:var(--gm3-sys-color-on-surface,#1f1f1f);opacity:0.38}.FAiUob .mIZh1c{background-color:var(--gm3-sys-color-outline,#747775)}.FAiUob .cXrdqd{background-color:#0b57d0;background-color:var(--gm3-sys-color-primary,#0b57d0)}.FAiUob .snByac{color:#444746;color:var(--gm3-sys-color-on-surface-variant,#444746)}.FAiUob.u3bW4e .snByac.snByac{color:#0b57d0;color:var(--gm3-sys-color-primary,#0b57d0)}.Em2Ord{margin:16px 0;outline:none}.Em2Ord+.Em2Ord{margin-top:24px}.Em2Ord:first-child{margin-top:0}.Em2Ord:last-child{margin-bottom:0}.PsAlOe{border-radius:8px;padding:16px}.PsAlOe>:first-child{margin-top:0}.PsAlOe>:last-child{margin-bottom:0}.PsAlOe .x9zgF{color:#1f1f1f;color:var(--gm3-sys-color-on-surface,#1f1f1f);font-family:"Google Sans",roboto,"Noto Sans Myanmar UI",arial,sans-serif;font-size:1rem;font-weight:500;letter-spacing:0rem;line-height:1.5}.PsAlOe.sj692e .x9zgF,.PsAlOe.sj692e .yTaH4c{color:#0842a0;color:var(--gm3-sys-color-on-primary-container,#0842a0)}.PsAlOe.Xq8bDe .x9zgF,.PsAlOe.Xq8bDe .yTaH4c{color:#410e0b;color:var(--gm3-sys-color-on-error-container,#8c1d18)}.PsAlOe.rNe0id .x9zgF,.PsAlOe.rNe0id .yTaH4c{color:var(--wf-color-warning-text,#421f00)}.PsAlOe .yTaH4c{color:#1f1f1f;color:var(--gm3-sys-color-on-surface,#1f1f1f)}.PsAlOe.YFdWic .vYeFie,.PsAlOe.YFdWic .yTaH4c{margin-left:64px;width:calc(100% - 48px - 16px)}.PsAlOe.YFdWic .yTaH4c{color:#444746;color:var(--gm3-sys-color-on-surface-variant,#444746);margin-top:4px}.PsAlOe.YFdWic:not(.S7S4N) .vYeFie{margin-left:0;width:0}.PsAlOe:not(.S7S4N)>.yTaH4c{margin-top:0}.PsAlOe.sj692e{background:#d3e3fd;background:var(--gm3-sys-color-primary-container,#d3e3fd)}.PsAlOe.Xq8bDe{background:#f9dedc;background:var(--gm3-sys-color-error-container,#f9dedc)}.PsAlOe.rNe0id{background:var(--wf-color-warning-bg,#fff0d1)}.PsAlOe.YFdWic{background:#f8fafd;background:var(--gm3-sys-color-surface-container-low,#f8fafd);min-height:80px;position:relative}.PsAlOe.YFdWic .x9zgF{color:#1f1f1f;color:var(--gm3-sys-color-on-surface,#1f1f1f)}.PsAlOe.YFdWic .yTaH4c{color:#444746;color:var(--gm3-sys-color-on-surface-variant,#444746)}.PsAlOe:not(.S7S4N){display:-webkit-box;display:-webkit-flex;display:flex}.Em2Ord.eLNT1d{display:none}.Em2Ord.RDPZE{opacity:.5;pointer-events:none}.Em2Ord.RDPZE .Em2Ord.RDPZE{opacity:1}.se0rCf{background-color:#f8fafd;background-color:var(--gm3-sys-color-surface-container-low,#f8fafd);border-radius:28px;padding:16px}.se0rCf .x9zgF{color:#1f1f1f;color:var(--gm3-sys-color-on-surface,#1f1f1f)}.se0rCf .yTaH4c{color:#444746;color:var(--gm3-sys-color-on-surface-variant,#444746)}.se0rCf .X3mtXb .snByac,.se0rCf.Em2Ord .i79UJc .snByac{background-color:#f8fafd;background-color:var(--gm3-sys-color-surface-container-low,#f8fafd)}.se0rCf .SgHwWb{display:-webkit-box;display:-webkit-flex;display:flex;-webkit-box-pack:end;-webkit-justify-content:flex-end;justify-content:flex-end;margin-top:16px}.se0rCf .SgHwWb .BqKGqe{margin-bottom:0;margin-top:0}.nn7x3d{border-bottom:1px solid #c4c7c5;border-bottom:1px solid var(--gm3-sys-color-outline-variant,#c4c7c5);display:-webkit-box;display:-webkit-flex;display:flex;-webkit-box-orient:vertical;-webkit-box-direction:normal;-webkit-flex-direction:column;flex-direction:column}.nn7x3d .V9RXW .rBUW7e{border-bottom:0}.nn7x3d .nn7x3d:last-child{border-bottom:0}.dwkQ3b:not(.jVwmLb){border-bottom:0}.nn7x3d .nn7x3d:last-child .ozEFYb{padding-bottom:0}.nn7x3d.dwkQ3b{border-bottom:0}.vYeFie:empty,.osxBFb:empty{display:none}.vYeFie>:first-child{margin-top:0;padding-top:0}.vYeFie>:last-child{margin-bottom:0;padding-bottom:0}.LwQQGe{margin:0 0 8px}.nn7x3d[data-expand-type="1"] .ozEFYb,.Em2Ord[data-expand-type="1"] .HKEKLe{cursor:pointer}.nn7x3d .ozEFYb{padding-bottom:16px}.x9zgF{-webkit-box-align:center;-webkit-align-items:center;align-items:center;color:#1f1f1f;color:var(--gm3-sys-color-on-surface,#1f1f1f);display:-webkit-box;display:-webkit-flex;display:flex;font-family:"Google Sans",roboto,"Noto Sans Myanmar UI",arial,sans-serif;font-size:1.25rem;font-weight:400;letter-spacing:0rem;line-height:1.2;margin-top:0;margin-bottom:0;padding:0}.Em2Ord.S7S4N .Em2Ord:not(.nn7x3d) .x9zgF{font-family:"Google Sans",roboto,"Noto Sans Myanmar UI",arial,sans-serif;font-size:1rem;font-weight:500;letter-spacing:0rem;line-height:1.5}.nn7x3d.u3bW4e .x9zgF{position:relative}.nn7x3d[data-expand-type="1"].u3bW4e .x9zgF::after{background:#0b57d0;background:var(--gm3-sys-color-primary,#0b57d0);border-radius:8px;bottom:-4px;content:"";left:-8px;position:absolute;opacity:0.1;right:-8px;top:-4px;z-index:-1}.HKEKLe{background:none;border:none;color:inherit;-webkit-box-flex:1;-webkit-flex-grow:1;flex-grow:1;font:inherit;margin:0;outline:0;padding:0;text-align:inherit}.HKEKLe::-moz-focus-inner{border:0}.HKEKLe [jsslot]{position:relative}.MI3XC{margin-left:16px}.MI3XC .aHWa4d{-webkit-box-align:center;-webkit-align-items:center;align-items:center;display:-webkit-box;display:-webkit-flex;display:flex;height:24px;-webkit-box-pack:center;-webkit-justify-content:center;justify-content:center;-webkit-transition:-webkit-transform 0.2s cubic-bezier(0.4,0,0.2,1);transition:-webkit-transform 0.2s cubic-bezier(0.4,0,0.2,1);transition:transform 0.2s cubic-bezier(0.4,0,0.2,1);transition:transform 0.2s cubic-bezier(0.4,0,0.2,1),-webkit-transform 0.2s cubic-bezier(0.4,0,0.2,1);width:24px}.nn7x3d .MI3XC,.nn7x3d .HKEKLe,.nn7x3d .CuWxc{pointer-events:none}.nn7x3d.jVwmLb .aHWa4d{-webkit-transform:rotate(-180deg);transform:rotate(-180deg)}.CuWxc{color:var(--gm3-sys-color-on-surface-variant,#444746);-webkit-flex-shrink:0;flex-shrink:0;height:20px;margin-right:16px;width:20px}.CuWxc .C3qbwe{height:100%;width:100%}.PsAlOe .CuWxc{margin-top:0}.PsAlOe.sj692e .CuWxc{color:#0b57d0;color:var(--gm3-sys-color-primary,#0b57d0)}.PsAlOe.Xq8bDe .CuWxc{color:#b3261e;color:var(--gm3-sys-color-error,#b3261e)}.PsAlOe.rNe0id .CuWxc{color:var(--wf-color-warning-icon,#f09d00)}.PsAlOe.YFdWic .CuWxc{height:48px;left:16px;position:absolute;top:16px;width:48px}.osxBFb{color:#444746;color:var(--gm3-sys-color-on-surface-variant,#444746);font-size:0.875rem;font-weight:400;line-height:1.4285714286;margin-top:8px}.vYeFie:empty+.yTaH4c{margin-top:0}.yTaH4c{margin-bottom:16px;margin-top:10px}.se0rCf .yTaH4c{margin-bottom:0;margin-top:16px}.yTaH4c:only-child{margin-bottom:0;margin-top:0}.nn7x3d .yTaH4c{margin-top:0;overflow:hidden;-webkit-transition:0.2s cubic-bezier(0.4,0,0.2,1);transition:0.2s cubic-bezier(0.4,0,0.2,1)}.nn7x3d.jVwmLb .yTaH4c{margin-bottom:0;margin-top:0;max-height:0;opacity:0;visibility:hidden}.yTaH4c>[jsslot]>:first-child:not(.PsAlOe){margin-top:0;padding-top:0}.yTaH4c>[jsslot]>:last-child:not(.PsAlOe){margin-bottom:0;padding-bottom:0}.kvM7xe{margin-bottom:-12px}.kvM7xe{-webkit-align-self:center;align-self:center;margin-bottom:0}.g0ndYb{border-bottom:1px solid #c4c7c5;border-bottom:1px solid var(--gm3-sys-color-outline-variant,#c4c7c5);display:-webkit-box;display:-webkit-flex;display:flex;-webkit-box-orient:horizontal;-webkit-box-direction:normal;-webkit-flex-direction:row;flex-direction:row;-webkit-box-pack:center;-webkit-justify-content:center;justify-content:center;height:0;margin-top:12px}.VXMllb{background-color:#fff;background-color:var(--gm3-sys-color-surface-container-lowest,#fff);display:-webkit-box;display:-webkit-flex;display:flex;height:24px;margin-top:-12px}.dwkQ3b:not(.jVwmLb) .g0ndYb{display:none}.dgtjld .VfPpkd-IE5DDf{background-color:#000;background-color:var(--gm3-sys-color-scrim,#000);opacity:0.32}.dgtjld .VfPpkd-P5QLlc{background-color:#e9eef6;background-color:var(--gm3-sys-color-surface-container-high,#e9eef6);border-radius:23px}.dgtjld .VfPpkd-k2Wrsb{color:#1f1f1f;color:var(--gm3-sys-color-on-surface,#1f1f1f);font-family:"Google Sans",roboto,"Noto Sans Myanmar UI",arial,sans-serif;font-size:1.5rem;font-weight:400;letter-spacing:0rem;line-height:1.3333333333}.dgtjld .VfPpkd-cnG4Wd{color:#444746;color:var(--gm3-sys-color-on-surface-variant,#444746);font-family:"Google Sans",roboto,"Noto Sans Myanmar UI",arial,sans-serif;font-size:0.875rem;font-weight:400;letter-spacing:0rem;line-height:1.4285714286;padding-bottom:0}.dgtjld .VfPpkd-T0kwCb{padding:0 24px 16px 24px}.dgtjld .yTaH4c{margin-left:0;margin-right:0;padding-left:0;padding-right:0}.dgtjld .ksBjEc.ksBjEc{color:#0b57d0;color:var(--gm3-sys-color-primary,#0b57d0);font-size:0.875rem;height:40px;padding:0 16px}.dgtjld .ksBjEc.ksBjEc:hover:not(:disabled){color:#0b57d0;color:var(--gm3-sys-color-primary,#0b57d0)}.dgtjld .ksBjEc.ksBjEc .VfPpkd-Jh9lGc::after,.dgtjld .ksBjEc.ksBjEc .VfPpkd-Jh9lGc::before{background-color:#0b57d0;background-color:var(--gm3-sys-color-primary,#0b57d0)}.dgtjld .ksBjEc.ksBjEc:focus:not(:disabled){color:#0b57d0;color:var(--gm3-sys-color-primary,#0b57d0)}.dgtjld .ksBjEc.ksBjEc .VfPpkd-J1Ukfc-LhBDec{border-color:#0b57d0;border-color:var(--gm3-sys-color-primary,#0b57d0)}.dgtjld .ksBjEc.ksBjEc .VfPpkd-J1Ukfc-LhBDec::after{border-color:#d3e3fd;border-color:var(--gm3-sys-color-primary-container,#d3e3fd)}.dgtjld .ksBjEc.ksBjEc .VfPpkd-J1Ukfc-LhBDec::after,.dgtjld .ksBjEc.ksBjEc .VfPpkd-J1Ukfc-LhBDec,.dgtjld .ksBjEc.ksBjEc .VfPpkd-Jh9lGc{border-radius:23px}.dgtjld.Zttm2{border-radius:0}.dgtjld.Zttm2 .VfPpkd-P5QLlc{height:100vh;max-height:none;max-width:none;width:100vw}.dgtjld.Zttm2 .yHy1rc{color:#444746;color:var(--gm3-sys-color-on-surface-variant,#444746);display:inline-block;padding:12px;text-align:center}.dgtjld.Zttm2 .VfPpkd-zMU9ub .NMm5M{fill:var(--gm3-sys-color-primary,#0b57d0)}.dgtjld.Zttm2 .VfPpkd-Bz112c-J1Ukfc-LhBDec{border-color:#0b57d0;border-color:var(--gm3-sys-color-primary,#0b57d0);padding:2px}.dgtjld.Zttm2 .VfPpkd-Bz112c-J1Ukfc-LhBDec,.dgtjld.Zttm2 .VfPpkd-Bz112c-J1Ukfc-LhBDec::after{border-radius:50%}.dgtjld.Zttm2 .yHy1rc:not(.VfPpkd-Bz112c-J1Ukfc-LhBDec)::before{display:none}.dgtjld.Zttm2 .yHy1rc:not(.VfPpkd-Bz112c-J1Ukfc-LhBDec)::after{background:none;border:none;box-shadow:none}.dgtjld.Zttm2 .yHy1rc .VfPpkd-Bz112c-Jh9lGc::before,.dgtjld.Zttm2 .yHy1rc .VfPpkd-Bz112c-Jh9lGc::after{background-color:#0b57d0;background-color:var(--gm3-sys-color-primary,#0b57d0)}.Zttm2 .rcN2gf{height:100%;width:100%}.Zttm2 .RITe7{border:none;color-scheme:normal;display:block;height:100%;padding:0;width:100%}.KGgLze{color:#444746;color:var(--gm3-sys-color-on-surface-variant,#444746);font-family:"Google Sans",roboto,"Noto Sans Myanmar UI",arial,sans-serif;-webkit-box-flex:1;-webkit-flex-grow:1;flex-grow:1;font-size:0.875rem;font-weight:400;padding-left:16px}.VfPpkd-JGcpL-uI4vCe-LkdAo,.VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:#6200ee;stroke:var(--mdc-theme-primary,#6200ee)}@media (-ms-high-contrast:active),screen and (forced-colors:active){.VfPpkd-JGcpL-uI4vCe-LkdAo,.VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:CanvasText}}.VfPpkd-JGcpL-uI4vCe-u014N{stroke:transparent}@-webkit-keyframes mdc-circular-progress-container-rotate{to{-webkit-transform:rotate(1turn);transform:rotate(1turn)}}@keyframes mdc-circular-progress-container-rotate{to{-webkit-transform:rotate(1turn);transform:rotate(1turn)}}@-webkit-keyframes mdc-circular-progress-spinner-layer-rotate{12.5%{-webkit-transform:rotate(135deg);transform:rotate(135deg)}25%{-webkit-transform:rotate(270deg);transform:rotate(270deg)}37.5%{-webkit-transform:rotate(405deg);transform:rotate(405deg)}50%{-webkit-transform:rotate(540deg);transform:rotate(540deg)}62.5%{-webkit-transform:rotate(675deg);transform:rotate(675deg)}75%{-webkit-transform:rotate(810deg);transform:rotate(810deg)}87.5%{-webkit-transform:rotate(945deg);transform:rotate(945deg)}100%{-webkit-transform:rotate(3turn);transform:rotate(3turn)}}@keyframes mdc-circular-progress-spinner-layer-rotate{12.5%{-webkit-transform:rotate(135deg);transform:rotate(135deg)}25%{-webkit-transform:rotate(270deg);transform:rotate(270deg)}37.5%{-webkit-transform:rotate(405deg);transform:rotate(405deg)}50%{-webkit-transform:rotate(540deg);transform:rotate(540deg)}62.5%{-webkit-transform:rotate(675deg);transform:rotate(675deg)}75%{-webkit-transform:rotate(810deg);transform:rotate(810deg)}87.5%{-webkit-transform:rotate(945deg);transform:rotate(945deg)}100%{-webkit-transform:rotate(3turn);transform:rotate(3turn)}}@-webkit-keyframes mdc-circular-progress-color-1-fade-in-out{from{opacity:.99}25%{opacity:.99}26%{opacity:0}89%{opacity:0}90%{opacity:.99}to{opacity:.99}}@keyframes mdc-circular-progress-color-1-fade-in-out{from{opacity:.99}25%{opacity:.99}26%{opacity:0}89%{opacity:0}90%{opacity:.99}to{opacity:.99}}@-webkit-keyframes mdc-circular-progress-color-2-fade-in-out{from{opacity:0}15%{opacity:0}25%{opacity:.99}50%{opacity:.99}51%{opacity:0}to{opacity:0}}@keyframes mdc-circular-progress-color-2-fade-in-out{from{opacity:0}15%{opacity:0}25%{opacity:.99}50%{opacity:.99}51%{opacity:0}to{opacity:0}}@-webkit-keyframes mdc-circular-progress-color-3-fade-in-out{from{opacity:0}40%{opacity:0}50%{opacity:.99}75%{opacity:.99}76%{opacity:0}to{opacity:0}}@keyframes mdc-circular-progress-color-3-fade-in-out{from{opacity:0}40%{opacity:0}50%{opacity:.99}75%{opacity:.99}76%{opacity:0}to{opacity:0}}@-webkit-keyframes mdc-circular-progress-color-4-fade-in-out{from{opacity:0}65%{opacity:0}75%{opacity:.99}90%{opacity:.99}to{opacity:0}}@keyframes mdc-circular-progress-color-4-fade-in-out{from{opacity:0}65%{opacity:0}75%{opacity:.99}90%{opacity:.99}to{opacity:0}}@-webkit-keyframes mdc-circular-progress-left-spin{from{-webkit-transform:rotate(265deg);transform:rotate(265deg)}50%{-webkit-transform:rotate(130deg);transform:rotate(130deg)}to{-webkit-transform:rotate(265deg);transform:rotate(265deg)}}@keyframes mdc-circular-progress-left-spin{from{-webkit-transform:rotate(265deg);transform:rotate(265deg)}50%{-webkit-transform:rotate(130deg);transform:rotate(130deg)}to{-webkit-transform:rotate(265deg);transform:rotate(265deg)}}@-webkit-keyframes mdc-circular-progress-right-spin{from{-webkit-transform:rotate(-265deg);transform:rotate(-265deg)}50%{-webkit-transform:rotate(-130deg);transform:rotate(-130deg)}to{-webkit-transform:rotate(-265deg);transform:rotate(-265deg)}}@keyframes mdc-circular-progress-right-spin{from{-webkit-transform:rotate(-265deg);transform:rotate(-265deg)}50%{-webkit-transform:rotate(-130deg);transform:rotate(-130deg)}to{-webkit-transform:rotate(-265deg);transform:rotate(-265deg)}}.VfPpkd-JGcpL-P1ekSe{display:-webkit-inline-box;display:-webkit-inline-flex;display:inline-flex;position:relative;direction:ltr;line-height:0;overflow:hidden;-webkit-transition:opacity .25s 0ms cubic-bezier(.4,0,.6,1);transition:opacity .25s 0ms cubic-bezier(.4,0,.6,1)}.VfPpkd-JGcpL-uI4vCe-haAclf,.VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G,.VfPpkd-JGcpL-IdXvz-haAclf,.VfPpkd-JGcpL-QYI5B-pbTTYe{position:absolute;width:100%;height:100%}.VfPpkd-JGcpL-uI4vCe-haAclf{-webkit-transform:rotate(-90deg);transform:rotate(-90deg)}.VfPpkd-JGcpL-IdXvz-haAclf{font-size:0;letter-spacing:0;white-space:nowrap;opacity:0}.VfPpkd-JGcpL-uI4vCe-LkdAo-Bd00G,.VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{fill:transparent}.VfPpkd-JGcpL-uI4vCe-LkdAo{-webkit-transition:stroke-dashoffset .5s 0ms cubic-bezier(0,0,.2,1);transition:stroke-dashoffset .5s 0ms cubic-bezier(0,0,.2,1)}.VfPpkd-JGcpL-OcUoKf-TpMipd{position:absolute;top:0;left:47.5%;box-sizing:border-box;width:5%;height:100%;overflow:hidden}.VfPpkd-JGcpL-OcUoKf-TpMipd .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{left:-900%;width:2000%;-webkit-transform:rotate(180deg);transform:rotate(180deg)}.VfPpkd-JGcpL-lLvYUc-e9ayKc{display:-webkit-inline-box;display:-webkit-inline-flex;display:inline-flex;position:relative;width:50%;height:100%;overflow:hidden}.VfPpkd-JGcpL-lLvYUc-e9ayKc .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{width:200%}.VfPpkd-JGcpL-lLvYUc-qwU8Me .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{left:-100%}.VfPpkd-JGcpL-P1ekSe-OWXEXe-A9y3zc .VfPpkd-JGcpL-uI4vCe-haAclf{opacity:0}.VfPpkd-JGcpL-P1ekSe-OWXEXe-A9y3zc .VfPpkd-JGcpL-IdXvz-haAclf{opacity:1}.VfPpkd-JGcpL-P1ekSe-OWXEXe-A9y3zc .VfPpkd-JGcpL-IdXvz-haAclf{-webkit-animation:mdc-circular-progress-container-rotate 1.5682352941176s linear infinite;animation:mdc-circular-progress-container-rotate 1.5682352941176s linear infinite}.VfPpkd-JGcpL-P1ekSe-OWXEXe-A9y3zc .VfPpkd-JGcpL-QYI5B-pbTTYe{-webkit-animation:mdc-circular-progress-spinner-layer-rotate 5332ms cubic-bezier(.4,0,.2,1) infinite both;animation:mdc-circular-progress-spinner-layer-rotate 5332ms cubic-bezier(.4,0,.2,1) infinite both}.VfPpkd-JGcpL-P1ekSe-OWXEXe-A9y3zc .VfPpkd-JGcpL-Ydhldb-R6PoUb{-webkit-animation:mdc-circular-progress-spinner-layer-rotate 5332ms cubic-bezier(.4,0,.2,1) infinite both,mdc-circular-progress-color-1-fade-in-out 5332ms cubic-bezier(.4,0,.2,1) infinite both;animation:mdc-circular-progress-spinner-layer-rotate 5332ms cubic-bezier(.4,0,.2,1) infinite both,mdc-circular-progress-color-1-fade-in-out 5332ms cubic-bezier(.4,0,.2,1) infinite both}.VfPpkd-JGcpL-P1ekSe-OWXEXe-A9y3zc .VfPpkd-JGcpL-Ydhldb-ibL1re{-webkit-animation:mdc-circular-progress-spinner-layer-rotate 5332ms cubic-bezier(.4,0,.2,1) infinite both,mdc-circular-progress-color-2-fade-in-out 5332ms cubic-bezier(.4,0,.2,1) infinite both;animation:mdc-circular-progress-spinner-layer-rotate 5332ms cubic-bezier(.4,0,.2,1) infinite both,mdc-circular-progress-color-2-fade-in-out 5332ms cubic-bezier(.4,0,.2,1) infinite both}.VfPpkd-JGcpL-P1ekSe-OWXEXe-A9y3zc .VfPpkd-JGcpL-Ydhldb-c5RTEf{-webkit-animation:mdc-circular-progress-spinner-layer-rotate 5332ms cubic-bezier(.4,0,.2,1) infinite both,mdc-circular-progress-color-3-fade-in-out 5332ms cubic-bezier(.4,0,.2,1) infinite both;animation:mdc-circular-progress-spinner-layer-rotate 5332ms cubic-bezier(.4,0,.2,1) infinite both,mdc-circular-progress-color-3-fade-in-out 5332ms cubic-bezier(.4,0,.2,1) infinite both}.VfPpkd-JGcpL-P1ekSe-OWXEXe-A9y3zc .VfPpkd-JGcpL-Ydhldb-II5mzb{-webkit-animation:mdc-circular-progress-spinner-layer-rotate 5332ms cubic-bezier(.4,0,.2,1) infinite both,mdc-circular-progress-color-4-fade-in-out 5332ms cubic-bezier(.4,0,.2,1) infinite both;animation:mdc-circular-progress-spinner-layer-rotate 5332ms cubic-bezier(.4,0,.2,1) infinite both,mdc-circular-progress-color-4-fade-in-out 5332ms cubic-bezier(.4,0,.2,1) infinite both}.VfPpkd-JGcpL-P1ekSe-OWXEXe-A9y3zc .VfPpkd-JGcpL-lLvYUc-LK5yu .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{-webkit-animation:mdc-circular-progress-left-spin 1333ms cubic-bezier(.4,0,.2,1) infinite both;animation:mdc-circular-progress-left-spin 1333ms cubic-bezier(.4,0,.2,1) infinite both}.VfPpkd-JGcpL-P1ekSe-OWXEXe-A9y3zc .VfPpkd-JGcpL-lLvYUc-qwU8Me .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{-webkit-animation:mdc-circular-progress-right-spin 1333ms cubic-bezier(.4,0,.2,1) infinite both;animation:mdc-circular-progress-right-spin 1333ms cubic-bezier(.4,0,.2,1) infinite both}.VfPpkd-JGcpL-P1ekSe-OWXEXe-xTMeO{opacity:0}.DU29of{position:relative}.DU29of .VfPpkd-JGcpL-uI4vCe-LkdAo,.DU29of .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:#4285f4}@media screen and (forced-colors:active),(-ms-high-contrast:active){.DU29of .VfPpkd-JGcpL-uI4vCe-LkdAo,.DU29of .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:CanvasText}}.DU29of .VfPpkd-JGcpL-Ydhldb-R6PoUb .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:#4285f4}@media screen and (forced-colors:active),(-ms-high-contrast:active){.DU29of .VfPpkd-JGcpL-Ydhldb-R6PoUb .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:CanvasText}}.DU29of .VfPpkd-JGcpL-Ydhldb-ibL1re .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:#ea4335}@media screen and (forced-colors:active),(-ms-high-contrast:active){.DU29of .VfPpkd-JGcpL-Ydhldb-ibL1re .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:CanvasText}}.DU29of .VfPpkd-JGcpL-Ydhldb-c5RTEf .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:#fbbc04}@media screen and (forced-colors:active),(-ms-high-contrast:active){.DU29of .VfPpkd-JGcpL-Ydhldb-c5RTEf .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:CanvasText}}.DU29of .VfPpkd-JGcpL-Ydhldb-II5mzb .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:#34a853}@media screen and (forced-colors:active),(-ms-high-contrast:active){.DU29of .VfPpkd-JGcpL-Ydhldb-II5mzb .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:CanvasText}}.DU29of .VfPpkd-JGcpL-Mr8B3-V67aGc{height:100%;width:100%;position:absolute;opacity:0;overflow:hidden;z-index:-1}.VfPpkd-BFbNVe-bF1uUb{position:absolute;border-radius:inherit;pointer-events:none;opacity:0;opacity:var(--mdc-elevation-overlay-opacity,0);-webkit-transition:opacity .28s cubic-bezier(.4,0,.2,1);transition:opacity .28s cubic-bezier(.4,0,.2,1);background-color:#fff;background-color:var(--mdc-elevation-overlay-color,#fff)}.NZp2ef{background-color:#e8eaed}.GY1Nfe{display:-webkit-inline-box;display:-webkit-inline-flex;display:inline-flex;place-content:center;place-items:center}html[dir=rtl] .giSqbe{-webkit-transform:scaleX(-1);transform:scaleX(-1)}.VfPpkd-z59Tgd{border-radius:4px;border-radius:var(--mdc-shape-small,4px)}.VfPpkd-Djsh7e-XxIAqe-ma6Yeb,.VfPpkd-Djsh7e-XxIAqe-cGMI2b{border-radius:4px;border-radius:var(--mdc-shape-small,4px)}.VfPpkd-z59Tgd{color:white;color:var(--mdc-theme-text-primary-on-dark,white)}.VfPpkd-z59Tgd{background-color:rgba(0,0,0,.6)}.VfPpkd-MlC99b{color:rgba(0,0,0,.87);color:var(--mdc-theme-text-primary-on-light,rgba(0,0,0,.87))}.VfPpkd-IqDDtd{color:rgba(0,0,0,.6)}.VfPpkd-IqDDtd-hSRGPd{color:#6200ee;color:var(--mdc-theme-primary,#6200ee)}.VfPpkd-a1tyJ-bN97Pc{overflow-x:unset;overflow-y:auto}.VfPpkd-suEOdc.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-z59Tgd,.VfPpkd-suEOdc.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-Djsh7e-XxIAqe-ma6Yeb,.VfPpkd-suEOdc.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-Djsh7e-XxIAqe-cGMI2b{background-color:#fff}.VfPpkd-z59Tgd{-moz-osx-font-smoothing:grayscale;-webkit-font-smoothing:antialiased;font-family:Roboto,sans-serif;font-family:var(--mdc-typography-caption-font-family,var(--mdc-typography-font-family,Roboto,sans-serif));font-size:.75rem;font-size:var(--mdc-typography-caption-font-size,.75rem);font-weight:400;font-weight:var(--mdc-typography-caption-font-weight,400);letter-spacing:.0333333333em;letter-spacing:var(--mdc-typography-caption-letter-spacing,.0333333333em);text-decoration:inherit;-webkit-text-decoration:var(--mdc-typography-caption-text-decoration,inherit);text-decoration:var(--mdc-typography-caption-text-decoration,inherit);text-transform:inherit;text-transform:var(--mdc-typography-caption-text-transform,inherit)}.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-z59Tgd{box-shadow:0 3px 1px -2px rgba(0,0,0,.2),0 2px 2px 0 rgba(0,0,0,.14),0 1px 5px 0 rgba(0,0,0,.12);border-radius:4px;line-height:20px}.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-z59Tgd .VfPpkd-BFbNVe-bF1uUb{width:100%;height:100%;top:0;left:0}.VfPpkd-z59Tgd .VfPpkd-MlC99b{display:block;margin-top:0;line-height:20px;-moz-osx-font-smoothing:grayscale;-webkit-font-smoothing:antialiased;font-family:Roboto,sans-serif;font-family:var(--mdc-typography-subtitle2-font-family,var(--mdc-typography-font-family,Roboto,sans-serif));font-size:.875rem;font-size:var(--mdc-typography-subtitle2-font-size,.875rem);line-height:1.375rem;line-height:var(--mdc-typography-subtitle2-line-height,1.375rem);font-weight:500;font-weight:var(--mdc-typography-subtitle2-font-weight,500);letter-spacing:.0071428571em;letter-spacing:var(--mdc-typography-subtitle2-letter-spacing,.0071428571em);text-decoration:inherit;-webkit-text-decoration:var(--mdc-typography-subtitle2-text-decoration,inherit);text-decoration:var(--mdc-typography-subtitle2-text-decoration,inherit);text-transform:inherit;text-transform:var(--mdc-typography-subtitle2-text-transform,inherit)}.VfPpkd-z59Tgd .VfPpkd-MlC99b::before{display:inline-block;width:0;height:24px;content:"";vertical-align:0}.VfPpkd-z59Tgd .VfPpkd-IqDDtd{-moz-osx-font-smoothing:grayscale;-webkit-font-smoothing:antialiased;font-family:Roboto,sans-serif;font-family:var(--mdc-typography-body2-font-family,var(--mdc-typography-font-family,Roboto,sans-serif));font-size:.875rem;font-size:var(--mdc-typography-body2-font-size,.875rem);line-height:1.25rem;line-height:var(--mdc-typography-body2-line-height,1.25rem);font-weight:400;font-weight:var(--mdc-typography-body2-font-weight,400);letter-spacing:.0178571429em;letter-spacing:var(--mdc-typography-body2-letter-spacing,.0178571429em);text-decoration:inherit;-webkit-text-decoration:var(--mdc-typography-body2-text-decoration,inherit);text-decoration:var(--mdc-typography-body2-text-decoration,inherit);text-transform:inherit;text-transform:var(--mdc-typography-body2-text-transform,inherit)}.VfPpkd-z59Tgd{word-break:break-all;word-break:var(--mdc-tooltip-word-break,normal);overflow-wrap:anywhere}.VfPpkd-suEOdc-OWXEXe-eo9XGd-RCfa3e .VfPpkd-z59Tgd-OiiCO{-webkit-transition:opacity .15s 0ms cubic-bezier(0,0,.2,1),-webkit-transform .15s 0ms cubic-bezier(0,0,.2,1);transition:opacity .15s 0ms cubic-bezier(0,0,.2,1),-webkit-transform .15s 0ms cubic-bezier(0,0,.2,1);transition:opacity .15s 0ms cubic-bezier(0,0,.2,1),transform .15s 0ms cubic-bezier(0,0,.2,1);transition:opacity .15s 0ms cubic-bezier(0,0,.2,1),transform .15s 0ms cubic-bezier(0,0,.2,1),-webkit-transform .15s 0ms cubic-bezier(0,0,.2,1)}.VfPpkd-suEOdc-OWXEXe-ZYIfFd-RCfa3e .VfPpkd-z59Tgd-OiiCO{-webkit-transition:opacity 75ms 0ms cubic-bezier(.4,0,1,1);transition:opacity 75ms 0ms cubic-bezier(.4,0,1,1)}.VfPpkd-suEOdc{position:fixed;display:none;z-index:9}.VfPpkd-suEOdc-sM5MNb-OWXEXe-nzrxxc{position:relative}.VfPpkd-suEOdc-OWXEXe-TSZdd,.VfPpkd-suEOdc-OWXEXe-eo9XGd,.VfPpkd-suEOdc-OWXEXe-ZYIfFd{display:-webkit-inline-box;display:-webkit-inline-flex;display:inline-flex}.VfPpkd-suEOdc-OWXEXe-TSZdd.VfPpkd-suEOdc-OWXEXe-nzrxxc,.VfPpkd-suEOdc-OWXEXe-eo9XGd.VfPpkd-suEOdc-OWXEXe-nzrxxc,.VfPpkd-suEOdc-OWXEXe-ZYIfFd.VfPpkd-suEOdc-OWXEXe-nzrxxc{display:inline-block;left:-320px;position:absolute}.VfPpkd-z59Tgd{line-height:16px;padding:4px 8px;min-width:40px;max-width:200px;min-height:24px;max-height:40vh;box-sizing:border-box;overflow:hidden;text-align:center}.VfPpkd-z59Tgd::before{position:absolute;box-sizing:border-box;width:100%;height:100%;top:0;left:0;border:1px solid transparent;border-radius:inherit;content:"";pointer-events:none}@media screen and (forced-colors:active){.VfPpkd-z59Tgd::before{border-color:CanvasText}}.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-z59Tgd{-webkit-box-align:start;-webkit-align-items:flex-start;align-items:flex-start;display:-webkit-box;display:-webkit-flex;display:flex;-webkit-box-orient:vertical;-webkit-box-direction:normal;-webkit-flex-direction:column;flex-direction:column;min-height:24px;min-width:40px;max-width:320px;position:relative;text-align:left}[dir=rtl] .VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-z59Tgd,.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-z59Tgd[dir=rtl]{text-align:right}.VfPpkd-suEOdc-OWXEXe-LlMNQd .VfPpkd-z59Tgd{text-align:left}[dir=rtl] .VfPpkd-suEOdc-OWXEXe-LlMNQd .VfPpkd-z59Tgd,.VfPpkd-suEOdc-OWXEXe-LlMNQd .VfPpkd-z59Tgd[dir=rtl]{text-align:right}.VfPpkd-z59Tgd .VfPpkd-MlC99b{margin:0 8px}.VfPpkd-z59Tgd .VfPpkd-IqDDtd{max-width:184px;margin:8px}.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-z59Tgd .VfPpkd-IqDDtd{max-width:304px;-webkit-align-self:stretch;align-self:stretch}.VfPpkd-z59Tgd .VfPpkd-IqDDtd-hSRGPd{text-decoration:none}.VfPpkd-suEOdc-OWXEXe-nzrxxc-LQLjdd,.VfPpkd-IqDDtd,.VfPpkd-MlC99b{z-index:1}.VfPpkd-z59Tgd-OiiCO{opacity:0;-webkit-transform:scale(.8);transform:scale(.8);will-change:transform,opacity}.VfPpkd-suEOdc-OWXEXe-TSZdd .VfPpkd-z59Tgd-OiiCO{-webkit-transform:scale(1);transform:scale(1);opacity:1}.VfPpkd-suEOdc-OWXEXe-ZYIfFd .VfPpkd-z59Tgd-OiiCO{-webkit-transform:scale(1);transform:scale(1)}.VfPpkd-Djsh7e-XxIAqe-ma6Yeb,.VfPpkd-Djsh7e-XxIAqe-cGMI2b{position:absolute;height:24px;width:24px;-webkit-transform:rotate(35deg) skewY(20deg) scaleX(.9396926208);transform:rotate(35deg) skewY(20deg) scaleX(.9396926208)}.VfPpkd-Djsh7e-XxIAqe-ma6Yeb .VfPpkd-BFbNVe-bF1uUb,.VfPpkd-Djsh7e-XxIAqe-cGMI2b .VfPpkd-BFbNVe-bF1uUb{width:100%;height:100%;top:0;left:0}.VfPpkd-Djsh7e-XxIAqe-cGMI2b{box-shadow:0 3px 1px -2px rgba(0,0,0,.2),0 2px 2px 0 rgba(0,0,0,.14),0 1px 5px 0 rgba(0,0,0,.12);outline:1px solid transparent;z-index:-1}@media screen and (forced-colors:active){.VfPpkd-Djsh7e-XxIAqe-cGMI2b{outline-color:CanvasText}}.EY8ABd{z-index:2101}.EY8ABd .VfPpkd-z59Tgd{background-color:#3c4043;color:#e8eaed}.EY8ABd .VfPpkd-MlC99b,.EY8ABd .VfPpkd-IqDDtd{color:#3c4043}.EY8ABd .VfPpkd-IqDDtd-hSRGPd{color:#1a73e8}.EY8ABd.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-z59Tgd,.EY8ABd.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-Djsh7e-XxIAqe-ma6Yeb,.EY8ABd.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-Djsh7e-XxIAqe-cGMI2b{background-color:#fff}.EY8ABd.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-MlC99b{font-family:"Google Sans",Roboto,Arial,sans-serif;line-height:1.25rem;font-size:.875rem;letter-spacing:.0178571429em;font-weight:500}.EY8ABd.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-z59Tgd{-webkit-border-radius:8px;border-radius:8px}.ziykHb{z-index:2101}.ziykHb .VfPpkd-z59Tgd{background-color:#3c4043;color:#e8eaed}.ziykHb .VfPpkd-MlC99b,.ziykHb .VfPpkd-IqDDtd{color:#3c4043}.ziykHb .VfPpkd-IqDDtd-hSRGPd{color:#1a73e8}.ziykHb.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-z59Tgd,.ziykHb.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-Djsh7e-XxIAqe-ma6Yeb,.ziykHb.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-Djsh7e-XxIAqe-cGMI2b{background-color:#fff}.ziykHb.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-MlC99b{font-family:"Google Sans",Roboto,Arial,sans-serif;line-height:1.25rem;font-size:.875rem;letter-spacing:.0178571429em;font-weight:500}.ziykHb.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-z59Tgd{-webkit-border-radius:8px;border-radius:8px}.EY8ABd-OWXEXe-TAWMXe{position:absolute;left:-10000px;top:auto;width:1px;height:1px;overflow:hidden;-webkit-user-select:none;-webkit-user-select:none}.NMm5M{fill:currentColor;-webkit-flex-shrink:0;flex-shrink:0}[dir=rtl] .hhikbc{-webkit-transform:scaleX(-1);transform:scaleX(-1)}.PrDSKc,.v42QC{padding-bottom:3px;padding-top:9px}.v42QC{margin:0}.PrDSKc:empty,.v42QC:empty{display:none}.TyDcZc,.jC5pMd{padding-bottom:3px;padding-top:9px}.jC5pMd{margin:0}.TyDcZc:empty,.jC5pMd:empty{display:none}.SXdXAb-BFbNVe,.SXdXAb-ugnUJb,.SXdXAb-BFbNVe::before,.SXdXAb-BFbNVe::after{border-radius:inherit;inset:0;position:absolute;pointer-events:none}.SXdXAb-ugnUJb{-webkit-transition:75ms opacity linear;transition:75ms opacity linear;background-color:var(--gm3-elevation-surface-tint-layer-color,transparent);opacity:calc(clamp(0, var(--gm3-elevation-level, 0), .05) + clamp(0, var(--gm3-elevation-level, 0) - 1, .03) + clamp(0, var(--gm3-elevation-level, 0) - 2, .03) + clamp(0, var(--gm3-elevation-level, 0) - 3, .01) + clamp(0, var(--gm3-elevation-level, 0) - 4, .02))}.SXdXAb-BFbNVe::before,.SXdXAb-BFbNVe::after{-webkit-transition:75ms box-shadow linear;transition:75ms box-shadow linear;content:""}.SXdXAb-BFbNVe::before{box-shadow:0 calc(1px*(clamp(0, var(--gm3-elevation-level, 0), 1) + clamp(0, var(--gm3-elevation-level, 0) - 3, 1) + clamp(0, var(--gm3-elevation-level, 0) - 4, 1)*2)) calc(1px*(2*clamp(0, var(--gm3-elevation-level, 0), 1) + clamp(0, var(--gm3-elevation-level, 0) - 2, 1) + clamp(0, var(--gm3-elevation-level, 0) - 4, 1))) 0 var(--gm3-elevation-shadow-color,transparent);opacity:calc(clamp(0, var(--gm3-elevation-level, 0), 1)*.3)}.SXdXAb-BFbNVe::after{box-shadow:0 calc(1px*(clamp(0, var(--gm3-elevation-level, 0), 1) + clamp(0, var(--gm3-elevation-level, 0) - 1, 1) + clamp(0, var(--gm3-elevation-level, 0) - 2, 3)*2)) calc(1px*(clamp(0, var(--gm3-elevation-level, 0), 2)*3 + clamp(0, var(--gm3-elevation-level, 0) - 2, 3)*2)) calc(1px*(clamp(0, var(--gm3-elevation-level, 0), 4) + 2*clamp(0, var(--gm3-elevation-level, 0) - 4, 1))) var(--gm3-elevation-shadow-color,transparent);opacity:calc(clamp(0, var(--gm3-elevation-level, 0), 1)*.15)}@media (forced-colors:active){.SXdXAb-BFbNVe{display:none}}.OiePBf-zPjgPe{display:var(--gm3-focus-ring-outward-display,none);pointer-events:none;position:absolute;z-index:1;border-start-start-radius:calc(var(--gm3-focus-ring-outward-target-shape-start-start, 0px) + var(--gm3-focus-ring-outward-offset, 2px));border-start-end-radius:calc(var(--gm3-focus-ring-outward-target-shape-start-end, 0px) + var(--gm3-focus-ring-outward-offset, 2px));border-end-end-radius:calc(var(--gm3-focus-ring-outward-target-shape-end-end, 0px) + var(--gm3-focus-ring-outward-offset, 2px));border-end-start-radius:calc(var(--gm3-focus-ring-outward-target-shape-end-start, 0px) + var(--gm3-focus-ring-outward-offset, 2px));inset:calc(var(--gm3-focus-ring-outward-offset, 2px)*-1);box-shadow:0 0 0 var(--gm3-focus-ring-outward-track-width,3px) var(--gm3-focus-ring-outward-color,var(--gm3-sys-color-secondary,#00639b));outline:var(--gm3-focus-ring-outward-track-width,3px) solid transparent;-webkit-animation-name:gm3-focus-ring-outward-grows,gm3-focus-ring-outward-shrinks;animation-name:gm3-focus-ring-outward-grows,gm3-focus-ring-outward-shrinks;-webkit-animation-duration:.15s,.45s;animation-duration:.15s,.45s;-webkit-animation-delay:0s,.15s;animation-delay:0s,.15s;-webkit-animation-timing-function:cubic-bezier(.2,0,0,1),cubic-bezier(.2,0,0,1);animation-timing-function:cubic-bezier(.2,0,0,1),cubic-bezier(.2,0,0,1)}@-webkit-keyframes gm3-focus-ring-outward-grows{from{box-shadow:0 0 0 0 var(--gm3-focus-ring-outward-color,var(--gm3-sys-color-secondary,#00639b))}to{box-shadow:0 0 0 8px var(--gm3-focus-ring-outward-color,var(--gm3-sys-color-secondary,#00639b))}}@keyframes gm3-focus-ring-outward-grows{from{box-shadow:0 0 0 0 var(--gm3-focus-ring-outward-color,var(--gm3-sys-color-secondary,#00639b))}to{box-shadow:0 0 0 8px var(--gm3-focus-ring-outward-color,var(--gm3-sys-color-secondary,#00639b))}}@-webkit-keyframes gm3-focus-ring-outward-shrinks{from{box-shadow:0 0 0 8px var(--gm3-focus-ring-outward-color,var(--gm3-sys-color-secondary,#00639b))}}@keyframes gm3-focus-ring-outward-shrinks{from{box-shadow:0 0 0 8px var(--gm3-focus-ring-outward-color,var(--gm3-sys-color-secondary,#00639b))}}@media (prefers-reduced-motion){.OiePBf-zPjgPe{-webkit-animation:none;animation:none}}.RBHQF-ksKsZd{overflow:hidden;outline:none;-webkit-tap-highlight-color:transparent}.RBHQF-ksKsZd,.RBHQF-ksKsZd::before,.RBHQF-ksKsZd::after{position:absolute;pointer-events:none;top:0;left:0;width:100%;height:100%;border-start-start-radius:var(--gm3-ripple-shape-start-start,inherit);border-start-end-radius:var(--gm3-ripple-shape-start-end,inherit);border-end-start-radius:var(--gm3-ripple-shape-end-start,inherit);border-end-end-radius:var(--gm3-ripple-shape-end-end,inherit)}.RBHQF-ksKsZd::before,.RBHQF-ksKsZd::after{opacity:0;content:""}.RBHQF-ksKsZd::before{-webkit-transition:opacity 75ms linear,border-radius var(--gm3-ripple-border-radius-transition-duration,0ms) linear;transition:opacity 75ms linear,border-radius var(--gm3-ripple-border-radius-transition-duration,0ms) linear;background-color:var(--gm3-ripple-hover-color,transparent)}.RBHQF-ksKsZd-OWXEXe-ZmdkE::before{opacity:var(--gm3-ripple-hover-opacity,0)}.RBHQF-ksKsZd::after{opacity:0;background:-webkit-radial-gradient(closest-side,var(--gm3-ripple-pressed-color,transparent) max(100% - 70px,65%),transparent 100%);background:radial-gradient(closest-side,var(--gm3-ripple-pressed-color,transparent) max(100% - 70px,65%),transparent 100%);-webkit-transition:opacity .25s linear,border-radius var(--gm3-ripple-border-radius-transition-duration,0ms) linear;transition:opacity .25s linear,border-radius var(--gm3-ripple-border-radius-transition-duration,0ms) linear;-webkit-transform-origin:center center;transform-origin:center center}.RBHQF-ksKsZd-OWXEXe-QDgCrf::after{-webkit-transition-duration:105ms;transition-duration:105ms;opacity:var(--gm3-ripple-pressed-opacity,0)}@media (forced-colors:active){.RBHQF-ksKsZd{display:none}}.UywwFc-LgbsSe{display:-webkit-inline-box;display:-webkit-inline-flex;display:inline-flex;position:relative;-webkit-box-align:center;-webkit-align-items:center;align-items:center;-webkit-box-pack:center;-webkit-justify-content:center;justify-content:center;box-sizing:border-box;border:none;outline:none;background:transparent;-webkit-appearance:none;appearance:none;line-height:inherit;text-rendering:inherit;-webkit-user-select:none;user-select:none;vertical-align:middle;cursor:pointer;min-inline-size:var(--gm3-button-filled-container-min-width,64px);padding-block:0;-webkit-padding-start:var(--gm3-button-filled-leading-space,24px);padding-inline-start:var(--gm3-button-filled-leading-space,24px);-webkit-padding-end:var(--gm3-button-filled-trailing-space,24px);padding-inline-end:var(--gm3-button-filled-trailing-space,24px);block-size:var(--gm3-button-filled-container-height,40px);border-radius:var(--gm3-button-filled-container-shape,9999px);--gm3-ripple-hover-color:var(--gm3-button-filled-hover-state-layer-color,var(--gm3-sys-color-on-primary,#fff));--gm3-ripple-hover-opacity:var(--gm3-button-filled-hover-state-layer-opacity,0.08);--gm3-ripple-pressed-color:var(--gm3-button-filled-hover-state-layer-color,var(--gm3-sys-color-on-primary,#fff));--gm3-ripple-pressed-opacity:var(--gm3-button-filled-pressed-state-layer-opacity,0.1);--gm3-focus-ring-outward-color:var(--gm3-button-filled-focus-indicator-color,var(--gm3-sys-color-secondary,#00639b));--gm3-focus-ring-outward-offset:var(--gm3-button-filled-focus-indicator-outline-offset,2px);--gm3-focus-ring-outward-track-width:var(--gm3-button-filled-focus-indicator-thickness,3px);--gm3-focus-ring-outward-target-shape-start-start:var(--gm3-button-filled-container-shape,9999px);--gm3-focus-ring-outward-target-shape-start-end:var(--gm3-button-filled-container-shape,9999px);--gm3-focus-ring-outward-target-shape-end-end:var(--gm3-button-filled-container-shape,9999px);--gm3-focus-ring-outward-target-shape-end-start:var(--gm3-button-filled-container-shape,9999px)}.UywwFc-mRLv6:focus-visible{outline:none}.UywwFc-LgbsSe:focus-visible,.UywwFc-mRLv6:focus-visible~.UywwFc-UHGRz{--gm3-focus-ring-outward-display:block}.UywwFc-LgbsSe:disabled{cursor:default;pointer-events:none;--gm3-ripple-hover-opacity:0;--gm3-ripple-pressed-opacity:0}.UywwFc-LgbsSe-OWXEXe-SfQLQb-suEOdc:disabled{pointer-events:auto}.UywwFc-LgbsSe[hidden]{display:none}.UywwFc-vQzf8d{position:relative;text-align:center;color:var(--gm3-button-filled-label-text-color,var(--gm3-sys-color-on-primary,#fff));font-size:var(--gm3-button-filled-label-text-size,.875rem);font-family:var(--gm3-button-filled-label-text-font,"Google Sans",Roboto,Arial,sans-serif);font-weight:var(--gm3-button-filled-label-text-weight,500);letter-spacing:var(--gm3-button-filled-label-text-tracking,0);-webkit-text-decoration:var(--gm3-button-filled-label-text-decoration,none);text-decoration:var(--gm3-button-filled-label-text-decoration,none);font-variation-settings:var(--gm3-button-filled-label-text-font-variation-settings,initial)}.UywwFc-kSE8rc-FoKg4d-sLO9V-YoZ4jf .UywwFc-vQzf8d{font-family:var(--gm3-button-filled-label-text-font,"Google Sans Flex","Google Sans Text","Google Sans",Roboto,Arial,sans-serif)}.UywwFc-LgbsSe:hover .UywwFc-vQzf8d{color:var(--gm3-button-filled-hover-label-text-color,var(--gm3-sys-color-on-primary,#fff))}.UywwFc-LgbsSe:focus-visible .UywwFc-vQzf8d{color:var(--gm3-button-filled-focus-label-text-color,var(--gm3-sys-color-on-primary,#fff))}.UywwFc-LgbsSe:active .UywwFc-vQzf8d{color:var(--gm3-button-filled-pressed-label-text-color,var(--gm3-sys-color-on-primary,#fff))}.UywwFc-LgbsSe:disabled .UywwFc-vQzf8d{color:var(--gm3-button-filled-disabled-label-text-color,rgba(var(--gm3-sys-color-on-surface-rgb,31,31,31),.38))}.UywwFc-LgbsSe-OWXEXe-zcdHbf .UywwFc-vQzf8d{white-space:nowrap;text-overflow:ellipsis;overflow:hidden}.UywwFc-LgbsSe-OWXEXe-Bz112c-M1Soyc{-webkit-padding-start:var(--gm3-button-filled-with-leading-icon-leading-space,16px);padding-inline-start:var(--gm3-button-filled-with-leading-icon-leading-space,16px);-webkit-padding-end:var(--gm3-button-filled-with-leading-icon-trailing-space,24px);padding-inline-end:var(--gm3-button-filled-with-leading-icon-trailing-space,24px)}.UywwFc-LgbsSe-OWXEXe-Bz112c-M1Soyc .UywwFc-kBDsod-Rtc0Jf i,.UywwFc-LgbsSe-OWXEXe-Bz112c-M1Soyc .UywwFc-kBDsod-Rtc0Jf img,.UywwFc-LgbsSe-OWXEXe-Bz112c-M1Soyc .UywwFc-kBDsod-Rtc0Jf svg{-webkit-margin-end:var(--gm3-button-filled-with-icon-icon-label-space,8px);margin-inline-end:var(--gm3-button-filled-with-icon-icon-label-space,8px)}.UywwFc-LgbsSe-OWXEXe-Bz112c-UbuQg{-webkit-padding-start:var(--gm3-button-filled-with-trailing-icon-leading-space,24px);padding-inline-start:var(--gm3-button-filled-with-trailing-icon-leading-space,24px);-webkit-padding-end:var(--gm3-button-filled-with-trailing-icon-trailing-space,16px);padding-inline-end:var(--gm3-button-filled-with-trailing-icon-trailing-space,16px)}.UywwFc-LgbsSe-OWXEXe-Bz112c-UbuQg .UywwFc-kBDsod-Rtc0Jf i,.UywwFc-LgbsSe-OWXEXe-Bz112c-UbuQg .UywwFc-kBDsod-Rtc0Jf img,.UywwFc-LgbsSe-OWXEXe-Bz112c-UbuQg .UywwFc-kBDsod-Rtc0Jf svg{-webkit-margin-start:var(--gm3-button-filled-with-icon-icon-label-space,8px);margin-inline-start:var(--gm3-button-filled-with-icon-icon-label-space,8px)}.UywwFc-kBDsod-Rtc0Jf{display:none;position:relative;line-height:0;color:var(--gm3-button-filled-with-icon-icon-color,var(--gm3-sys-color-on-primary,#fff))}.UywwFc-kBDsod-Rtc0Jf i,.UywwFc-kBDsod-Rtc0Jf img,.UywwFc-kBDsod-Rtc0Jf svg{display:-webkit-inline-box;display:-webkit-inline-flex;display:inline-flex;position:relative;direction:inherit;color:inherit;font-size:var(--gm3-button-filled-with-icon-icon-size,18px);inline-size:var(--gm3-button-filled-with-icon-icon-size,18px);block-size:var(--gm3-button-filled-with-icon-icon-size,18px)}.UywwFc-LgbsSe:hover .UywwFc-kBDsod-Rtc0Jf{color:var(--gm3-button-filled-with-icon-hover-icon-color,var(--gm3-sys-color-on-primary,#fff))}.UywwFc-LgbsSe:focus-visible .UywwFc-kBDsod-Rtc0Jf{color:var(--gm3-button-filled-with-icon-focus-icon-color,var(--gm3-sys-color-on-primary,#fff))}.UywwFc-LgbsSe:active .UywwFc-kBDsod-Rtc0Jf{color:var(--gm3-button-filled-with-icon-pressed-icon-color,var(--gm3-sys-color-on-primary,#fff))}.UywwFc-LgbsSe:disabled .UywwFc-kBDsod-Rtc0Jf{color:var(--gm3-button-filled-with-icon-disabled-icon-color,rgba(var(--gm3-sys-color-on-surface-rgb,31,31,31),.38))}[dir=rtl] .UywwFc-LgbsSe-OWXEXe-drxrmf-Bz112c .UywwFc-kBDsod-Rtc0Jf,.UywwFc-LgbsSe-OWXEXe-drxrmf-Bz112c .UywwFc-kBDsod-Rtc0Jf[dir=rtl]{-webkit-transform:scaleX(-1);transform:scaleX(-1)}.UywwFc-LgbsSe-OWXEXe-Bz112c-M1Soyc .UywwFc-kBDsod-Rtc0Jf-OWXEXe-M1Soyc,.UywwFc-LgbsSe-OWXEXe-Bz112c-UbuQg .UywwFc-kBDsod-Rtc0Jf-OWXEXe-UbuQg{display:-webkit-inline-box;display:-webkit-inline-flex;display:inline-flex}.UywwFc-mRLv6{position:absolute;inset:0}.UywwFc-LgbsSe-OWXEXe-dgl2Hf{margin-block:max((48px - var(--gm3-button-filled-container-height,40px))/2,0px)}.UywwFc-RLmnJb{position:absolute;inline-size:max(48px,100%);block-size:max(48px,100%);inset:unset;top:50%;left:50%;-webkit-transform:translate(-50%,-50%);transform:translate(-50%,-50%)}.UywwFc-LgbsSe{will-change:transform,opacity;background-color:var(--gm3-button-filled-container-color,var(--gm3-sys-color-primary,#0b57d0));--gm3-elevation-level:var(--gm3-button-filled-container-elevation,0);--gm3-elevation-shadow-color:var(--gm3-button-filled-container-shadow-color,var(--gm3-sys-color-shadow,#000))}.UywwFc-LgbsSe:hover{--gm3-elevation-level:var(--gm3-button-filled-hover-container-elevation,1)}.UywwFc-LgbsSe:focus-visible{--gm3-elevation-level:var(--gm3-button-filled-focus-container-elevation,0)}.UywwFc-LgbsSe:active{--gm3-elevation-level:var(--gm3-button-filled-pressed-container-elevation,0)}.UywwFc-LgbsSe:disabled{background-color:var(--gm3-button-filled-disabled-container-color,rgba(var(--gm3-sys-color-on-surface-rgb,31,31,31),.12));--gm3-elevation-level:var(--gm3-button-filled-disabled-container-elevation,0)}.UywwFc-LgbsSe::before{content:"";pointer-events:none;position:absolute;inset:0;border-radius:inherit;border:1px solid transparent}@media (forced-colors:active){.UywwFc-LgbsSe:disabled::before{border-color:GrayText}}@media (forced-colors:active){.UywwFc-StrnGf-YYd4I-VtOx3e::before{border-color:CanvasText}}.ne2Ple-suEOdc{position:fixed;display:none;z-index:var(--gm3-tooltip-plain-z-index,2101)}.ne2Ple-z59Tgd{box-sizing:border-box;min-block-size:24px;min-inline-size:40px;overflow-wrap:anywhere;overflow:hidden;padding-block:4px;padding-inline:8px;word-break:normal;max-block-size:var(--gm3-tooltip-plain-container-max-block-size,40vh)}.ne2Ple-z59Tgd::before{position:absolute;box-sizing:border-box;inline-size:100%;block-size:100%;inset-block-start:0;inset-inline-start:0;border:1px solid transparent;border-radius:inherit;content:"";pointer-events:none}.ne2Ple-suEOdc-OWXEXe-TSZdd,.ne2Ple-suEOdc-OWXEXe-eo9XGd,.ne2Ple-suEOdc-OWXEXe-ZYIfFd{display:-webkit-inline-box;display:-webkit-inline-flex;display:inline-flex}.ne2Ple-z59Tgd-OiiCO{opacity:0;-webkit-transform:scale(.8);transform:scale(.8);will-change:transform,opacity}.ne2Ple-suEOdc-OWXEXe-TSZdd .ne2Ple-z59Tgd-OiiCO{opacity:1;-webkit-transform:scale(1);transform:scale(1)}.ne2Ple-suEOdc-OWXEXe-ZYIfFd .ne2Ple-z59Tgd-OiiCO{-webkit-transform:scale(1);transform:scale(1)}.ne2Ple-suEOdc-OWXEXe-eo9XGd-RCfa3e .ne2Ple-z59Tgd-OiiCO{-webkit-transition:opacity .15s 0ms cubic-bezier(0,0,.2,1),-webkit-transform .15s 0ms cubic-bezier(0,0,.2,1);transition:opacity .15s 0ms cubic-bezier(0,0,.2,1),-webkit-transform .15s 0ms cubic-bezier(0,0,.2,1);transition:opacity .15s 0ms cubic-bezier(0,0,.2,1),transform .15s 0ms cubic-bezier(0,0,.2,1);transition:opacity .15s 0ms cubic-bezier(0,0,.2,1),transform .15s 0ms cubic-bezier(0,0,.2,1),-webkit-transform .15s 0ms cubic-bezier(0,0,.2,1)}.ne2Ple-suEOdc-OWXEXe-ZYIfFd-RCfa3e .ne2Ple-z59Tgd-OiiCO{-webkit-transition:opacity 75ms 0ms cubic-bezier(.4,0,1,1);transition:opacity 75ms 0ms cubic-bezier(.4,0,1,1)}.ne2Ple-suEOdc-OWXEXe-pijamc .ne2Ple-z59Tgd{max-inline-size:200px;background-color:var(--gm3-tooltip-plain-container-color,var(--gm3-sys-color-inverse-surface,#303030));border-radius:var(--gm3-tooltip-plain-container-shape,4px);color:var(--gm3-tooltip-plain-supporting-text-color,var(--gm3-sys-color-inverse-on-surface,#f2f2f2));font-family:var(--gm3-tooltip-plain-supporting-text-font,"Google Sans Text","Google Sans");font-size:var(--gm3-tooltip-plain-supporting-text-size,.75rem);font-weight:var(--gm3-tooltip-plain-supporting-text-weight,400);letter-spacing:var(--gm3-tooltip-plain-supporting-text-tracking,.00625rem);line-height:var(--gm3-tooltip-plain-supporting-text-line-height,1rem);text-align:center}.ne2Ple-suEOdc-OWXEXe-LlMNQd .ne2Ple-z59Tgd{text-align:start}.ne2Ple-oshW8e-V67aGc{position:absolute;left:-10000px;top:auto;inline-size:1px;height:1px;overflow:hidden;-webkit-user-select:none;user-select:none}.AeBiU-LgbsSe{display:-webkit-inline-box;display:-webkit-inline-flex;display:inline-flex;position:relative;-webkit-box-align:center;-webkit-align-items:center;align-items:center;-webkit-box-pack:center;-webkit-justify-content:center;justify-content:center;box-sizing:border-box;border:none;outline:none;background:transparent;-webkit-appearance:none;appearance:none;line-height:inherit;text-rendering:inherit;-webkit-user-select:none;user-select:none;vertical-align:middle;cursor:pointer;min-inline-size:var(--gm3-button-outlined-container-min-width,64px);padding-block:0;-webkit-padding-start:var(--gm3-button-outlined-leading-space,24px);padding-inline-start:var(--gm3-button-outlined-leading-space,24px);-webkit-padding-end:var(--gm3-button-outlined-trailing-space,24px);padding-inline-end:var(--gm3-button-outlined-trailing-space,24px);block-size:var(--gm3-button-outlined-container-height,40px);border-radius:var(--gm3-button-outlined-container-shape,9999px);--gm3-ripple-hover-color:var(--gm3-button-outlined-hover-state-layer-color,var(--gm3-sys-color-primary,#0b57d0));--gm3-ripple-hover-opacity:var(--gm3-button-outlined-hover-state-layer-opacity,0.08);--gm3-ripple-pressed-color:var(--gm3-button-outlined-hover-state-layer-color,var(--gm3-sys-color-primary,#0b57d0));--gm3-ripple-pressed-opacity:var(--gm3-button-outlined-pressed-state-layer-opacity,0.1);--gm3-focus-ring-outward-color:var(--gm3-button-outlined-focus-indicator-color,var(--gm3-sys-color-secondary,#00639b));--gm3-focus-ring-outward-offset:var(--gm3-button-outlined-focus-indicator-outline-offset,2px);--gm3-focus-ring-outward-track-width:var(--gm3-button-outlined-focus-indicator-thickness,3px);--gm3-focus-ring-outward-target-shape-start-start:var(--gm3-button-outlined-container-shape,9999px);--gm3-focus-ring-outward-target-shape-start-end:var(--gm3-button-outlined-container-shape,9999px);--gm3-focus-ring-outward-target-shape-end-end:var(--gm3-button-outlined-container-shape,9999px);--gm3-focus-ring-outward-target-shape-end-start:var(--gm3-button-outlined-container-shape,9999px)}.AeBiU-mRLv6:focus-visible{outline:none}.AeBiU-LgbsSe:focus-visible,.AeBiU-mRLv6:focus-visible~.AeBiU-UHGRz{--gm3-focus-ring-outward-display:block}.AeBiU-LgbsSe:disabled{cursor:default;pointer-events:none;--gm3-ripple-hover-opacity:0;--gm3-ripple-pressed-opacity:0}.AeBiU-LgbsSe-OWXEXe-SfQLQb-suEOdc:disabled{pointer-events:auto}.AeBiU-LgbsSe[hidden]{display:none}.AeBiU-vQzf8d{position:relative;text-align:center;color:var(--gm3-button-outlined-label-text-color,var(--gm3-sys-color-primary,#0b57d0));font-size:var(--gm3-button-outlined-label-text-size,.875rem);font-family:var(--gm3-button-outlined-label-text-font,"Google Sans",Roboto,Arial,sans-serif);font-weight:var(--gm3-button-outlined-label-text-weight,500);letter-spacing:var(--gm3-button-outlined-label-text-tracking,0);-webkit-text-decoration:var(--gm3-button-outlined-label-text-decoration,none);text-decoration:var(--gm3-button-outlined-label-text-decoration,none);font-variation-settings:var(--gm3-button-outlined-label-text-font-variation-settings,initial)}.AeBiU-kSE8rc-FoKg4d-sLO9V-YoZ4jf .AeBiU-vQzf8d{font-family:var(--gm3-button-outlined-label-text-font,"Google Sans Flex","Google Sans Text","Google Sans",Roboto,Arial,sans-serif)}.AeBiU-LgbsSe:hover .AeBiU-vQzf8d{color:var(--gm3-button-outlined-hover-label-text-color,var(--gm3-sys-color-primary,#0b57d0))}.AeBiU-LgbsSe:focus-visible .AeBiU-vQzf8d{color:var(--gm3-button-outlined-focus-label-text-color,var(--gm3-sys-color-primary,#0b57d0))}.AeBiU-LgbsSe:active .AeBiU-vQzf8d{color:var(--gm3-button-outlined-pressed-label-text-color,var(--gm3-sys-color-primary,#0b57d0))}.AeBiU-LgbsSe:disabled .AeBiU-vQzf8d{color:var(--gm3-button-outlined-disabled-label-text-color,rgba(var(--gm3-sys-color-on-surface-rgb,31,31,31),.38))}.AeBiU-LgbsSe-OWXEXe-zcdHbf .AeBiU-vQzf8d{white-space:nowrap;text-overflow:ellipsis;overflow:hidden}.AeBiU-LgbsSe-OWXEXe-Bz112c-M1Soyc{-webkit-padding-start:var(--gm3-button-outlined-with-leading-icon-leading-space,16px);padding-inline-start:var(--gm3-button-outlined-with-leading-icon-leading-space,16px);-webkit-padding-end:var(--gm3-button-outlined-with-leading-icon-trailing-space,24px);padding-inline-end:var(--gm3-button-outlined-with-leading-icon-trailing-space,24px)}.AeBiU-LgbsSe-OWXEXe-Bz112c-M1Soyc .AeBiU-kBDsod-Rtc0Jf i,.AeBiU-LgbsSe-OWXEXe-Bz112c-M1Soyc .AeBiU-kBDsod-Rtc0Jf img,.AeBiU-LgbsSe-OWXEXe-Bz112c-M1Soyc .AeBiU-kBDsod-Rtc0Jf svg{-webkit-margin-end:var(--gm3-button-outlined-with-icon-icon-label-space,8px);margin-inline-end:var(--gm3-button-outlined-with-icon-icon-label-space,8px)}.AeBiU-LgbsSe-OWXEXe-Bz112c-UbuQg{-webkit-padding-start:var(--gm3-button-outlined-with-trailing-icon-leading-space,24px);padding-inline-start:var(--gm3-button-outlined-with-trailing-icon-leading-space,24px);-webkit-padding-end:var(--gm3-button-outlined-with-trailing-icon-trailing-space,16px);padding-inline-end:var(--gm3-button-outlined-with-trailing-icon-trailing-space,16px)}.AeBiU-LgbsSe-OWXEXe-Bz112c-UbuQg .AeBiU-kBDsod-Rtc0Jf i,.AeBiU-LgbsSe-OWXEXe-Bz112c-UbuQg .AeBiU-kBDsod-Rtc0Jf img,.AeBiU-LgbsSe-OWXEXe-Bz112c-UbuQg .AeBiU-kBDsod-Rtc0Jf svg{-webkit-margin-start:var(--gm3-button-outlined-with-icon-icon-label-space,8px);margin-inline-start:var(--gm3-button-outlined-with-icon-icon-label-space,8px)}.AeBiU-kBDsod-Rtc0Jf{display:none;position:relative;line-height:0;color:var(--gm3-button-outlined-with-icon-icon-color,var(--gm3-sys-color-primary,#0b57d0))}.AeBiU-kBDsod-Rtc0Jf i,.AeBiU-kBDsod-Rtc0Jf img,.AeBiU-kBDsod-Rtc0Jf svg{display:-webkit-inline-box;display:-webkit-inline-flex;display:inline-flex;position:relative;direction:inherit;color:inherit;font-size:var(--gm3-button-outlined-with-icon-icon-size,18px);inline-size:var(--gm3-button-outlined-with-icon-icon-size,18px);block-size:var(--gm3-button-outlined-with-icon-icon-size,18px)}.AeBiU-LgbsSe:hover .AeBiU-kBDsod-Rtc0Jf{color:var(--gm3-button-outlined-with-icon-hover-icon-color,var(--gm3-sys-color-primary,#0b57d0))}.AeBiU-LgbsSe:focus-visible .AeBiU-kBDsod-Rtc0Jf{color:var(--gm3-button-outlined-with-icon-focus-icon-color,var(--gm3-sys-color-primary,#0b57d0))}.AeBiU-LgbsSe:active .AeBiU-kBDsod-Rtc0Jf{color:var(--gm3-button-outlined-with-icon-pressed-icon-color,var(--gm3-sys-color-primary,#0b57d0))}.AeBiU-LgbsSe:disabled .AeBiU-kBDsod-Rtc0Jf{color:var(--gm3-button-outlined-with-icon-disabled-icon-color,rgba(var(--gm3-sys-color-on-surface-rgb,31,31,31),.38))}[dir=rtl] .AeBiU-LgbsSe-OWXEXe-drxrmf-Bz112c .AeBiU-kBDsod-Rtc0Jf,.AeBiU-LgbsSe-OWXEXe-drxrmf-Bz112c .AeBiU-kBDsod-Rtc0Jf[dir=rtl]{-webkit-transform:scaleX(-1);transform:scaleX(-1)}.AeBiU-LgbsSe-OWXEXe-Bz112c-M1Soyc .AeBiU-kBDsod-Rtc0Jf-OWXEXe-M1Soyc,.AeBiU-LgbsSe-OWXEXe-Bz112c-UbuQg .AeBiU-kBDsod-Rtc0Jf-OWXEXe-UbuQg{display:-webkit-inline-box;display:-webkit-inline-flex;display:inline-flex}.AeBiU-mRLv6{position:absolute;inset:0}.AeBiU-LgbsSe-OWXEXe-dgl2Hf{margin-block:max((48px - var(--gm3-button-outlined-container-height,40px))/2,0px)}.AeBiU-RLmnJb{position:absolute;inline-size:max(48px,100%);block-size:max(48px,100%);inset:unset;top:50%;left:50%;-webkit-transform:translate(-50%,-50%);transform:translate(-50%,-50%)}.AeBiU-LgbsSe{border-style:solid;border-width:var(--gm3-button-outlined-outline-width,1px);border-color:var(--gm3-button-outlined-outline-color,var(--gm3-sys-color-outline,#747775));--gm3-focus-ring-outward-offset:calc(var(--gm3-button-outlined-focus-indicator-outline-offset, 2px) + var(--gm3-button-outlined-outline-width, 1px));--gm3-focus-ring-outward-target-shape-start-start:calc(var(--gm3-button-outlined-container-shape, 9999px) - var(--gm3-button-outlined-outline-width, 1px));--gm3-focus-ring-outward-target-shape-start-end:calc(var(--gm3-button-outlined-container-shape, 9999px) - var(--gm3-button-outlined-outline-width, 1px));--gm3-focus-ring-outward-target-shape-end-end:calc(var(--gm3-button-outlined-container-shape, 9999px) - var(--gm3-button-outlined-outline-width, 1px));--gm3-focus-ring-outward-target-shape-end-start:calc(var(--gm3-button-outlined-container-shape, 9999px) - var(--gm3-button-outlined-outline-width, 1px))}.AeBiU-LgbsSe:hover{border-color:var(--gm3-button-outlined-hover-outline-color,var(--gm3-sys-color-outline,#747775))}.AeBiU-LgbsSe:focus-visible{border-color:var(--gm3-button-outlined-focus-outline-color,var(--gm3-sys-color-primary,#0b57d0))}.AeBiU-LgbsSe:active{border-color:var(--gm3-button-outlined-pressed-outline-color,var(--gm3-sys-color-outline,#747775))}.AeBiU-LgbsSe:disabled{border-color:var(--gm3-button-outlined-disabled-outline-color,rgba(var(--gm3-sys-color-on-surface-rgb,31,31,31),.12))}@media (forced-colors:active){.AeBiU-LgbsSe:disabled{border-color:GrayText}}.AeBiU-RLmnJb{inline-size:max(48px,100% + var(--gm3-button-outlined-outline-width,1px) * 2)}.mUIrbf-LgbsSe{display:-webkit-inline-box;display:-webkit-inline-flex;display:inline-flex;position:relative;-webkit-box-align:center;-webkit-align-items:center;align-items:center;-webkit-box-pack:center;-webkit-justify-content:center;justify-content:center;box-sizing:border-box;border:none;outline:none;background:transparent;-webkit-appearance:none;appearance:none;line-height:inherit;text-rendering:inherit;-webkit-user-select:none;user-select:none;vertical-align:middle;cursor:pointer;min-inline-size:var(--gm3-button-text-container-min-width,64px);padding-block:0;-webkit-padding-start:var(--gm3-button-text-leading-space,12px);padding-inline-start:var(--gm3-button-text-leading-space,12px);-webkit-padding-end:var(--gm3-button-text-trailing-space,12px);padding-inline-end:var(--gm3-button-text-trailing-space,12px);block-size:var(--gm3-button-text-container-height,40px);border-radius:var(--gm3-button-text-container-shape,9999px);--gm3-ripple-hover-color:var(--gm3-button-text-hover-state-layer-color,var(--gm3-sys-color-primary,#0b57d0));--gm3-ripple-hover-opacity:var(--gm3-button-text-hover-state-layer-opacity,0.08);--gm3-ripple-pressed-color:var(--gm3-button-text-hover-state-layer-color,var(--gm3-sys-color-primary,#0b57d0));--gm3-ripple-pressed-opacity:var(--gm3-button-text-pressed-state-layer-opacity,0.1);--gm3-focus-ring-outward-color:var(--gm3-button-text-focus-indicator-color,var(--gm3-sys-color-secondary,#00639b));--gm3-focus-ring-outward-offset:var(--gm3-button-text-focus-indicator-outline-offset,2px);--gm3-focus-ring-outward-track-width:var(--gm3-button-text-focus-indicator-thickness,3px);--gm3-focus-ring-outward-target-shape-start-start:var(--gm3-button-text-container-shape,9999px);--gm3-focus-ring-outward-target-shape-start-end:var(--gm3-button-text-container-shape,9999px);--gm3-focus-ring-outward-target-shape-end-end:var(--gm3-button-text-container-shape,9999px);--gm3-focus-ring-outward-target-shape-end-start:var(--gm3-button-text-container-shape,9999px)}.mUIrbf-mRLv6:focus-visible{outline:none}.mUIrbf-LgbsSe:focus-visible,.mUIrbf-mRLv6:focus-visible~.mUIrbf-UHGRz{--gm3-focus-ring-outward-display:block}.mUIrbf-LgbsSe:disabled{cursor:default;pointer-events:none;--gm3-ripple-hover-opacity:0;--gm3-ripple-pressed-opacity:0}.mUIrbf-LgbsSe-OWXEXe-SfQLQb-suEOdc:disabled{pointer-events:auto}.mUIrbf-LgbsSe[hidden]{display:none}.mUIrbf-vQzf8d{position:relative;text-align:center;color:var(--gm3-button-text-label-text-color,var(--gm3-sys-color-primary,#0b57d0));font-size:var(--gm3-button-text-label-text-size,.875rem);font-family:var(--gm3-button-text-label-text-font,"Google Sans",Roboto,Arial,sans-serif);font-weight:var(--gm3-button-text-label-text-weight,500);letter-spacing:var(--gm3-button-text-label-text-tracking,0);-webkit-text-decoration:var(--gm3-button-text-label-text-decoration,none);text-decoration:var(--gm3-button-text-label-text-decoration,none);font-variation-settings:var(--gm3-button-text-label-text-font-variation-settings,initial)}.mUIrbf-kSE8rc-FoKg4d-sLO9V-YoZ4jf .mUIrbf-vQzf8d{font-family:var(--gm3-button-text-label-text-font,"Google Sans Flex","Google Sans Text","Google Sans",Roboto,Arial,sans-serif)}.mUIrbf-LgbsSe:hover .mUIrbf-vQzf8d{color:var(--gm3-button-text-hover-label-text-color,var(--gm3-sys-color-primary,#0b57d0))}.mUIrbf-LgbsSe:focus-visible .mUIrbf-vQzf8d{color:var(--gm3-button-text-focus-label-text-color,var(--gm3-sys-color-primary,#0b57d0))}.mUIrbf-LgbsSe:active .mUIrbf-vQzf8d{color:var(--gm3-button-text-pressed-label-text-color,var(--gm3-sys-color-primary,#0b57d0))}.mUIrbf-LgbsSe:disabled .mUIrbf-vQzf8d{color:var(--gm3-button-text-disabled-label-text-color,rgba(var(--gm3-sys-color-on-surface-rgb,31,31,31),.38))}.mUIrbf-LgbsSe-OWXEXe-zcdHbf .mUIrbf-vQzf8d{white-space:nowrap;text-overflow:ellipsis;overflow:hidden}.mUIrbf-LgbsSe-OWXEXe-Bz112c-M1Soyc{-webkit-padding-start:var(--gm3-button-text-with-leading-icon-leading-space,12px);padding-inline-start:var(--gm3-button-text-with-leading-icon-leading-space,12px);-webkit-padding-end:var(--gm3-button-text-with-leading-icon-trailing-space,16px);padding-inline-end:var(--gm3-button-text-with-leading-icon-trailing-space,16px)}.mUIrbf-LgbsSe-OWXEXe-Bz112c-M1Soyc .mUIrbf-kBDsod-Rtc0Jf i,.mUIrbf-LgbsSe-OWXEXe-Bz112c-M1Soyc .mUIrbf-kBDsod-Rtc0Jf img,.mUIrbf-LgbsSe-OWXEXe-Bz112c-M1Soyc .mUIrbf-kBDsod-Rtc0Jf svg{-webkit-margin-end:var(--gm3-button-text-with-icon-icon-label-space,8px);margin-inline-end:var(--gm3-button-text-with-icon-icon-label-space,8px)}.mUIrbf-LgbsSe-OWXEXe-Bz112c-UbuQg{-webkit-padding-start:var(--gm3-button-text-with-trailing-icon-leading-space,16px);padding-inline-start:var(--gm3-button-text-with-trailing-icon-leading-space,16px);-webkit-padding-end:var(--gm3-button-text-with-trailing-icon-trailing-space,12px);padding-inline-end:var(--gm3-button-text-with-trailing-icon-trailing-space,12px)}.mUIrbf-LgbsSe-OWXEXe-Bz112c-UbuQg .mUIrbf-kBDsod-Rtc0Jf i,.mUIrbf-LgbsSe-OWXEXe-Bz112c-UbuQg .mUIrbf-kBDsod-Rtc0Jf img,.mUIrbf-LgbsSe-OWXEXe-Bz112c-UbuQg .mUIrbf-kBDsod-Rtc0Jf svg{-webkit-margin-start:var(--gm3-button-text-with-icon-icon-label-space,8px);margin-inline-start:var(--gm3-button-text-with-icon-icon-label-space,8px)}.mUIrbf-kBDsod-Rtc0Jf{display:none;position:relative;line-height:0;color:var(--gm3-button-text-with-icon-icon-color,var(--gm3-sys-color-primary,#0b57d0))}.mUIrbf-kBDsod-Rtc0Jf i,.mUIrbf-kBDsod-Rtc0Jf img,.mUIrbf-kBDsod-Rtc0Jf svg{display:-webkit-inline-box;display:-webkit-inline-flex;display:inline-flex;position:relative;direction:inherit;color:inherit;font-size:var(--gm3-button-text-with-icon-icon-size,18px);inline-size:var(--gm3-button-text-with-icon-icon-size,18px);block-size:var(--gm3-button-text-with-icon-icon-size,18px)}.mUIrbf-LgbsSe:hover .mUIrbf-kBDsod-Rtc0Jf{color:var(--gm3-button-text-with-icon-hover-icon-color,var(--gm3-sys-color-primary,#0b57d0))}.mUIrbf-LgbsSe:focus-visible .mUIrbf-kBDsod-Rtc0Jf{color:var(--gm3-button-text-with-icon-focus-icon-color,var(--gm3-sys-color-primary,#0b57d0))}.mUIrbf-LgbsSe:active .mUIrbf-kBDsod-Rtc0Jf{color:var(--gm3-button-text-with-icon-pressed-icon-color,var(--gm3-sys-color-primary,#0b57d0))}.mUIrbf-LgbsSe:disabled .mUIrbf-kBDsod-Rtc0Jf{color:var(--gm3-button-text-with-icon-disabled-icon-color,rgba(var(--gm3-sys-color-on-surface-rgb,31,31,31),.38))}[dir=rtl] .mUIrbf-LgbsSe-OWXEXe-drxrmf-Bz112c .mUIrbf-kBDsod-Rtc0Jf,.mUIrbf-LgbsSe-OWXEXe-drxrmf-Bz112c .mUIrbf-kBDsod-Rtc0Jf[dir=rtl]{-webkit-transform:scaleX(-1);transform:scaleX(-1)}.mUIrbf-LgbsSe-OWXEXe-Bz112c-M1Soyc .mUIrbf-kBDsod-Rtc0Jf-OWXEXe-M1Soyc,.mUIrbf-LgbsSe-OWXEXe-Bz112c-UbuQg .mUIrbf-kBDsod-Rtc0Jf-OWXEXe-UbuQg{display:-webkit-inline-box;display:-webkit-inline-flex;display:inline-flex}.mUIrbf-mRLv6{position:absolute;inset:0}.mUIrbf-LgbsSe-OWXEXe-dgl2Hf{margin-block:max((48px - var(--gm3-button-text-container-height,40px))/2,0px)}.mUIrbf-RLmnJb{position:absolute;inline-size:max(48px,100%);block-size:max(48px,100%);inset:unset;top:50%;left:50%;-webkit-transform:translate(-50%,-50%);transform:translate(-50%,-50%)}.mUIrbf-LgbsSe{will-change:transform,opacity}.mUIrbf-LgbsSe::before{content:"";pointer-events:none;position:absolute;inset:0;border-radius:inherit;border:1px solid transparent}@media (forced-colors:active){.mUIrbf-LgbsSe:disabled::before{border-color:GrayText}}@media (forced-colors:active){.mUIrbf-StrnGf-YYd4I-VtOx3e::before{border-color:CanvasText}}.FOBRw-LgbsSe{display:-webkit-inline-box;display:-webkit-inline-flex;display:inline-flex;position:relative;-webkit-box-align:center;-webkit-align-items:center;align-items:center;-webkit-box-pack:center;-webkit-justify-content:center;justify-content:center;box-sizing:border-box;border:none;outline:none;background:transparent;-webkit-appearance:none;appearance:none;line-height:inherit;text-rendering:inherit;-webkit-user-select:none;user-select:none;vertical-align:middle;cursor:pointer;min-inline-size:var(--gm3-button-filled-tonal-container-min-width,64px);padding-block:0;-webkit-padding-start:var(--gm3-button-filled-tonal-leading-space,24px);padding-inline-start:var(--gm3-button-filled-tonal-leading-space,24px);-webkit-padding-end:var(--gm3-button-filled-tonal-trailing-space,24px);padding-inline-end:var(--gm3-button-filled-tonal-trailing-space,24px);block-size:var(--gm3-button-filled-tonal-container-height,40px);border-radius:var(--gm3-button-filled-tonal-container-shape,9999px);--gm3-ripple-hover-color:var(--gm3-button-filled-tonal-hover-state-layer-color,var(--gm3-sys-color-on-secondary-container,#001d35));--gm3-ripple-hover-opacity:var(--gm3-button-filled-tonal-hover-state-layer-opacity,0.08);--gm3-ripple-pressed-color:var(--gm3-button-filled-tonal-hover-state-layer-color,var(--gm3-sys-color-on-secondary-container,#001d35));--gm3-ripple-pressed-opacity:var(--gm3-button-filled-tonal-pressed-state-layer-opacity,0.1);--gm3-focus-ring-outward-color:var(--gm3-button-filled-tonal-focus-indicator-color,var(--gm3-sys-color-secondary,#00639b));--gm3-focus-ring-outward-offset:var(--gm3-button-filled-tonal-focus-indicator-outline-offset,2px);--gm3-focus-ring-outward-track-width:var(--gm3-button-filled-tonal-focus-indicator-thickness,3px);--gm3-focus-ring-outward-target-shape-start-start:var(--gm3-button-filled-tonal-container-shape,9999px);--gm3-focus-ring-outward-target-shape-start-end:var(--gm3-button-filled-tonal-container-shape,9999px);--gm3-focus-ring-outward-target-shape-end-end:var(--gm3-button-filled-tonal-container-shape,9999px);--gm3-focus-ring-outward-target-shape-end-start:var(--gm3-button-filled-tonal-container-shape,9999px)}.FOBRw-mRLv6:focus-visible{outline:none}.FOBRw-LgbsSe:focus-visible,.FOBRw-mRLv6:focus-visible~.FOBRw-UHGRz{--gm3-focus-ring-outward-display:block}.FOBRw-LgbsSe:disabled{cursor:default;pointer-events:none;--gm3-ripple-hover-opacity:0;--gm3-ripple-pressed-opacity:0}.FOBRw-LgbsSe-OWXEXe-SfQLQb-suEOdc:disabled{pointer-events:auto}.FOBRw-LgbsSe[hidden]{display:none}.FOBRw-vQzf8d{position:relative;text-align:center;color:var(--gm3-button-filled-tonal-label-text-color,var(--gm3-sys-color-on-secondary-container,#001d35));font-size:var(--gm3-button-filled-tonal-label-text-size,.875rem);font-family:var(--gm3-button-filled-tonal-label-text-font,"Google Sans",Roboto,Arial,sans-serif);font-weight:var(--gm3-button-filled-tonal-label-text-weight,500);letter-spacing:var(--gm3-button-filled-tonal-label-text-tracking,0);-webkit-text-decoration:var(--gm3-button-filled-tonal-label-text-decoration,none);text-decoration:var(--gm3-button-filled-tonal-label-text-decoration,none);font-variation-settings:var(--gm3-button-filled-tonal-label-text-font-variation-settings,initial)}.FOBRw-kSE8rc-FoKg4d-sLO9V-YoZ4jf .FOBRw-vQzf8d{font-family:var(--gm3-button-filled-tonal-label-text-font,"Google Sans Flex","Google Sans Text","Google Sans",Roboto,Arial,sans-serif)}.FOBRw-LgbsSe:hover .FOBRw-vQzf8d{color:var(--gm3-button-filled-tonal-hover-label-text-color,var(--gm3-sys-color-on-secondary-container,#001d35))}.FOBRw-LgbsSe:focus-visible .FOBRw-vQzf8d{color:var(--gm3-button-filled-tonal-focus-label-text-color,var(--gm3-sys-color-on-secondary-container,#001d35))}.FOBRw-LgbsSe:active .FOBRw-vQzf8d{color:var(--gm3-button-filled-tonal-pressed-label-text-color,var(--gm3-sys-color-on-secondary-container,#001d35))}.FOBRw-LgbsSe:disabled .FOBRw-vQzf8d{color:var(--gm3-button-filled-tonal-disabled-label-text-color,rgba(var(--gm3-sys-color-on-surface-rgb,31,31,31),.38))}.FOBRw-LgbsSe-OWXEXe-zcdHbf .FOBRw-vQzf8d{white-space:nowrap;text-overflow:ellipsis;overflow:hidden}.FOBRw-LgbsSe-OWXEXe-Bz112c-M1Soyc{-webkit-padding-start:var(--gm3-button-filled-tonal-with-leading-icon-leading-space,16px);padding-inline-start:var(--gm3-button-filled-tonal-with-leading-icon-leading-space,16px);-webkit-padding-end:var(--gm3-button-filled-tonal-with-leading-icon-trailing-space,24px);padding-inline-end:var(--gm3-button-filled-tonal-with-leading-icon-trailing-space,24px)}.FOBRw-LgbsSe-OWXEXe-Bz112c-M1Soyc .FOBRw-kBDsod-Rtc0Jf i,.FOBRw-LgbsSe-OWXEXe-Bz112c-M1Soyc .FOBRw-kBDsod-Rtc0Jf img,.FOBRw-LgbsSe-OWXEXe-Bz112c-M1Soyc .FOBRw-kBDsod-Rtc0Jf svg{-webkit-margin-end:var(--gm3-button-filled-tonal-with-icon-icon-label-space,8px);margin-inline-end:var(--gm3-button-filled-tonal-with-icon-icon-label-space,8px)}.FOBRw-LgbsSe-OWXEXe-Bz112c-UbuQg{-webkit-padding-start:var(--gm3-button-filled-tonal-with-trailing-icon-leading-space,24px);padding-inline-start:var(--gm3-button-filled-tonal-with-trailing-icon-leading-space,24px);-webkit-padding-end:var(--gm3-button-filled-tonal-with-trailing-icon-trailing-space,16px);padding-inline-end:var(--gm3-button-filled-tonal-with-trailing-icon-trailing-space,16px)}.FOBRw-LgbsSe-OWXEXe-Bz112c-UbuQg .FOBRw-kBDsod-Rtc0Jf i,.FOBRw-LgbsSe-OWXEXe-Bz112c-UbuQg .FOBRw-kBDsod-Rtc0Jf img,.FOBRw-LgbsSe-OWXEXe-Bz112c-UbuQg .FOBRw-kBDsod-Rtc0Jf svg{-webkit-margin-start:var(--gm3-button-filled-tonal-with-icon-icon-label-space,8px);margin-inline-start:var(--gm3-button-filled-tonal-with-icon-icon-label-space,8px)}.FOBRw-kBDsod-Rtc0Jf{display:none;position:relative;line-height:0;color:var(--gm3-button-filled-tonal-with-icon-icon-color,var(--gm3-sys-color-on-secondary-container,#001d35))}.FOBRw-kBDsod-Rtc0Jf i,.FOBRw-kBDsod-Rtc0Jf img,.FOBRw-kBDsod-Rtc0Jf svg{display:-webkit-inline-box;display:-webkit-inline-flex;display:inline-flex;position:relative;direction:inherit;color:inherit;font-size:var(--gm3-button-filled-tonal-with-icon-icon-size,18px);inline-size:var(--gm3-button-filled-tonal-with-icon-icon-size,18px);block-size:var(--gm3-button-filled-tonal-with-icon-icon-size,18px)}.FOBRw-LgbsSe:hover .FOBRw-kBDsod-Rtc0Jf{color:var(--gm3-button-filled-tonal-with-icon-hover-icon-color,var(--gm3-sys-color-on-secondary-container,#001d35))}.FOBRw-LgbsSe:focus-visible .FOBRw-kBDsod-Rtc0Jf{color:var(--gm3-button-filled-tonal-with-icon-focus-icon-color,var(--gm3-sys-color-on-secondary-container,#001d35))}.FOBRw-LgbsSe:active .FOBRw-kBDsod-Rtc0Jf{color:var(--gm3-button-filled-tonal-with-icon-pressed-icon-color,var(--gm3-sys-color-on-secondary-container,#001d35))}.FOBRw-LgbsSe:disabled .FOBRw-kBDsod-Rtc0Jf{color:var(--gm3-button-filled-tonal-with-icon-disabled-icon-color,rgba(var(--gm3-sys-color-on-surface-rgb,31,31,31),.38))}[dir=rtl] .FOBRw-LgbsSe-OWXEXe-drxrmf-Bz112c .FOBRw-kBDsod-Rtc0Jf,.FOBRw-LgbsSe-OWXEXe-drxrmf-Bz112c .FOBRw-kBDsod-Rtc0Jf[dir=rtl]{-webkit-transform:scaleX(-1);transform:scaleX(-1)}.FOBRw-LgbsSe-OWXEXe-Bz112c-M1Soyc .FOBRw-kBDsod-Rtc0Jf-OWXEXe-M1Soyc,.FOBRw-LgbsSe-OWXEXe-Bz112c-UbuQg .FOBRw-kBDsod-Rtc0Jf-OWXEXe-UbuQg{display:-webkit-inline-box;display:-webkit-inline-flex;display:inline-flex}.FOBRw-mRLv6{position:absolute;inset:0}.FOBRw-LgbsSe-OWXEXe-dgl2Hf{margin-block:max((48px - var(--gm3-button-filled-tonal-container-height,40px))/2,0px)}.FOBRw-RLmnJb{position:absolute;inline-size:max(48px,100%);block-size:max(48px,100%);inset:unset;top:50%;left:50%;-webkit-transform:translate(-50%,-50%);transform:translate(-50%,-50%)}.FOBRw-LgbsSe{will-change:transform,opacity;background-color:var(--gm3-button-filled-tonal-container-color,var(--gm3-sys-color-secondary-container,#c2e7ff));--gm3-elevation-level:var(--gm3-button-filled-tonal-container-elevation,0);--gm3-elevation-shadow-color:var(--gm3-button-filled-tonal-container-shadow-color,var(--gm3-sys-color-shadow,#000))}.FOBRw-LgbsSe:hover{--gm3-elevation-level:var(--gm3-button-filled-tonal-hover-container-elevation,1)}.FOBRw-LgbsSe:focus-visible{--gm3-elevation-level:var(--gm3-button-filled-tonal-focus-container-elevation,0)}.FOBRw-LgbsSe:active{--gm3-elevation-level:var(--gm3-button-filled-tonal-pressed-container-elevation,0)}.FOBRw-LgbsSe:disabled{background-color:var(--gm3-button-filled-tonal-disabled-container-color,rgba(var(--gm3-sys-color-on-surface-rgb,31,31,31),.12));--gm3-elevation-level:var(--gm3-button-filled-tonal-disabled-container-elevation,0)}.FOBRw-LgbsSe::before{content:"";pointer-events:none;position:absolute;inset:0;border-radius:inherit;border:1px solid transparent}@media (forced-colors:active){.FOBRw-LgbsSe:disabled::before{border-color:GrayText}}@media (forced-colors:active){.FOBRw-StrnGf-YYd4I-VtOx3e::before{border-color:CanvasText}}.tB5Jxf-xl07Ob-XxIAqe{display:none;position:absolute;box-sizing:border-box;margin:0;padding:0;border-radius:4px;-webkit-transform:scale(1);transform:scale(1);-webkit-transform-origin:top left;transform-origin:top left;opacity:0;will-change:transform,opacity;-webkit-transition:opacity .03s linear,height .25s cubic-bezier(0,0,.2,1),-webkit-transform .12s cubic-bezier(0,0,.2,1);transition:opacity .03s linear,height .25s cubic-bezier(0,0,.2,1),-webkit-transform .12s cubic-bezier(0,0,.2,1);transition:opacity .03s linear,transform .12s cubic-bezier(0,0,.2,1),height .25s cubic-bezier(0,0,.2,1);transition:opacity .03s linear,transform .12s cubic-bezier(0,0,.2,1),height .25s cubic-bezier(0,0,.2,1),-webkit-transform .12s cubic-bezier(0,0,.2,1);z-index:8;--gm3-elevation-level:var(--gm3-menu-surface-container-elevation,2);--gm3-elevation-shadow-color:var(--gm3-menu-surface-container-shadow-color,var(--gm3-sys-color-shadow,#000));max-width:calc(100vw - 32px);max-height:calc(100vw - 32px);background-color:var(--gm3-menu-surface-container-color,var(--gm3-sys-color-surface-container,#f0f4f9));color:#000}[dir=rtl] .tB5Jxf-xl07Ob-XxIAqe,.tB5Jxf-xl07Ob-XxIAqe[dir=rtl]{-webkit-transform-origin:top right;transform-origin:top right}.tB5Jxf-xl07Ob-XxIAqe-OWXEXe-Vkfede-QBLLGd{width:100%}.tB5Jxf-xl07Ob-S5Cmsd{overflow:auto;max-height:inherit;border-radius:inherit}.tB5Jxf-xl07Ob-XxIAqe:focus{outline:none}.tB5Jxf-xl07Ob-XxIAqe-OWXEXe-oT9UPb-FNFY6c{display:inline-block;-webkit-transform:scale(.8);transform:scale(.8);opacity:0}.tB5Jxf-xl07Ob-XxIAqe-OWXEXe-FNFY6c{display:inline-block;-webkit-transform:scale(1);transform:scale(1);opacity:1}.tB5Jxf-xl07Ob-XxIAqe-OWXEXe-oT9UPb-xTMeO{display:inline-block;opacity:0;-webkit-transition:opacity 75ms linear;transition:opacity 75ms linear}.tB5Jxf-xl07Ob-XxIAqe-OWXEXe-oYxtQd{position:relative;overflow:visible}.tB5Jxf-xl07Ob-XxIAqe-OWXEXe-qbOKL{position:fixed}.tB5Jxf-xl07Ob-XxIAqe-OWXEXe-uxVfW-FNFY6c-uFfGwd{border-start-start-radius:0;border-start-end-radius:0}.dMNVAe,.FSdAW{padding-bottom:3px;padding-top:9px}.FSdAW{margin:0}.dMNVAe:empty,.FSdAW:empty{display:none}@media screen and (prefers-color-scheme:dark){:root{--wf-color-warning-bg:#754200;--wf-color-warning-icon:#ffdf99;--wf-color-warning-text:#fff0d1}}@media screen and (prefers-color-scheme:light){:root{--wf-color-warning-bg:#fff0d1;--wf-color-warning-icon:#f09d00;--wf-color-warning-text:#421f00}}.hZUije{border:0}.hZUije.WS4XDd{max-height:1.3333em;padding:0 2px;vertical-align:middle;width:auto}.kHluYc{border:0;object-fit:contain}.kHluYc.WS4XDd{max-height:1.3333em;padding:0 2px;vertical-align:middle;width:auto}.vOZun,.gomQac{padding-bottom:3px;padding-top:9px;margin-bottom:0;margin-top:0}.gomQac{margin:0}.vOZun:empty{display:none}.JnOM6e{background-color:transparent;border:none;border-radius:4px;box-sizing:border-box;display:inline-block;font-size:14px;height:36px;letter-spacing:.15px;line-height:34px;padding:0 24px;position:relative;text-align:center}.JnOM6e:focus-visible{outline:none;position:relative}.JnOM6e:focus-visible::after{border:2px solid rgb(24,90,188);border-radius:6px;bottom:-4px;box-shadow:0 0 0 2px rgb(232,240,254);content:"";left:-4px;position:absolute;right:-4px;top:-4px}.rDisVe:focus:not(:focus-visible),.GjFdVe:focus:not(:focus-visible){box-shadow:0 1px 1px 0 rgba(66,133,244,.3),0 1px 3px 1px rgba(66,133,244,.15)}.rDisVe:hover:not(:focus-visible),.GjFdVe:hover:not(:focus-visible){box-shadow:0 1px 1px 0 rgba(66,133,244,.45),0 1px 3px 1px rgba(66,133,244,.3)}.JnOM6e:disabled{pointer-events:none}.JnOM6e:hover{cursor:pointer}.JnOM6e.kTeh9{line-height:36px;text-decoration:none}.JnOM6e.eLNT1d{display:none}.rDisVe{background-color:rgb(26,115,232);color:#fff}.rDisVe:disabled{background-color:rgb(232,234,237);color:rgb(154,160,166)}.rDisVe:focus,.rDisVe:hover{background-color:rgb(24,90,188)}.GjFdVe{border:1px solid rgb(218,220,224);color:rgb(26,115,232)}.GjFdVe:disabled{color:rgb(189,193,198)}.GjFdVe:active{background-color:rgb(174,203,250);color:rgb(23,78,166)}.GjFdVe:focus{background-color:rgb(232,240,254);border-color:rgb(24,90,188);color:rgb(23,78,166)}.GjFdVe:hover{background-color:rgb(232,240,254);color:rgb(23,78,166)}.KXbQ4b{color:rgb(26,115,232);min-width:0;padding-left:8px;padding-right:8px}.KXbQ4b:disabled{color:rgb(189,193,198)}.KXbQ4b:active,.KXbQ4b:hover{color:rgb(24,90,188)}.KXbQ4b:active{background-color:rgba(26,115,232,.12)}.KXbQ4b:focus,.KXbQ4b:hover{background-color:rgba(26,115,232,.04)}.aN1Vld{margin:16px 0;outline:none}.aN1Vld+.aN1Vld{margin-top:24px}.aN1Vld:first-child{margin-top:0}.aN1Vld:last-child{margin-bottom:0}.fegW5d{border-radius:8px;padding:16px}.fegW5d>:first-child{margin-top:0}.fegW5d>:last-child{margin-bottom:0}.fegW5d .cySqRb,.fegW5d .yOnVIb{color:rgb(32,33,36)}.fegW5d.YFdWic .yOnVIb{color:rgb(95,99,104);margin-top:4px;padding:0}.fegW5d.YFdWic .wSQNd,.fegW5d.YFdWic .yOnVIb{margin-left:64px;width:calc(100% - 64px)}.fegW5d.YFdWic:not(.S7S4N) .wSQNd{margin-left:0;width:0}.fegW5d:not(.S7S4N)>.yOnVIb{margin-top:0}.fegW5d.sj692e{background:rgb(232,240,254)}.fegW5d.Xq8bDe{background:rgb(252,232,230)}.fegW5d.rNe0id{background:rgb(254,247,224)}.fegW5d.YFdWic{border:1px solid rgb(218,220,224);min-height:80px;position:relative}.fegW5d:not(.S7S4N){display:-webkit-box;display:-webkit-flex;display:flex}.aN1Vld.eLNT1d{display:none}.aN1Vld.RDPZE{opacity:.5;pointer-events:none}.aN1Vld.RDPZE .aN1Vld.RDPZE{opacity:1}.wlrzMe{border:1px solid rgb(218,220,224);border-radius:8px;padding:16px}.wlrzMe .EEiyWe{display:-webkit-box;display:-webkit-flex;display:flex;-webkit-box-pack:end;-webkit-justify-content:flex-end;justify-content:flex-end;margin-top:16px}.wlrzMe .EEiyWe .GjFdVe{margin-bottom:0;margin-top:0}.wSQNd:empty{display:none}.wSQNd>:first-child{margin-top:0;padding-top:0}.wSQNd>:last-child{margin-bottom:0;padding-bottom:0}.cySqRb{-webkit-box-align:center;-webkit-align-items:center;align-items:center;color:rgb(32,33,36);display:-webkit-box;display:-webkit-flex;display:flex;font-size:16px;font-weight:500;letter-spacing:.1px;line-height:1.4286;margin-bottom:0;margin-top:0;padding:0}.zlrrr{color:rgb(95,99,104);-webkit-flex-shrink:0;flex-shrink:0;height:20px;margin-right:16px;width:20px}.zlrrr .GxLRef{height:100%;width:100%}.fegW5d .zlrrr{margin-top:0}.fegW5d.sj692e .zlrrr{color:rgb(25,103,210)}.fegW5d.Xq8bDe .zlrrr{color:rgb(197,34,31)}.fegW5d.rNe0id .zlrrr{color:rgb(234,134,0)}.fegW5d.YFdWic .zlrrr{height:48px;left:16px;position:absolute;top:16px;width:48px}.yOnVIb{margin:auto -24px;padding-left:24px;padding-right:24px;margin-bottom:16px;margin-top:10px}.wlrzMe .yOnVIb{margin-bottom:0;margin-top:16px}.yOnVIb>:first-child:not(section){margin-top:0;padding-top:0}.yOnVIb>:last-child:not(section){margin-bottom:0;padding-bottom:0}.wSQNd:empty+.yOnVIb{margin-top:0}.yOnVIb:only-child{margin-bottom:0;margin-top:0}c-wiz{contain:style}c-wiz>c-data{display:none}c-wiz.rETSD{contain:none}c-wiz.Ubi8Z{contain:layout style}.llhEMd{-webkit-transition:opacity .15s cubic-bezier(0.4,0,0.2,1) .15s;transition:opacity .15s cubic-bezier(0.4,0,0.2,1) .15s;background-color:rgba(0,0,0,0.502);bottom:0;left:0;opacity:0;position:fixed;right:0;top:0;z-index:5000}.llhEMd.iWO5td{-webkit-transition:opacity .05s cubic-bezier(0.4,0,0.2,1);transition:opacity .05s cubic-bezier(0.4,0,0.2,1);opacity:1}.mjANdc{transition:-webkit-transform .4s cubic-bezier(0.4,0,0.2,1);-webkit-transition:-webkit-transform .4s cubic-bezier(0.4,0,0.2,1);-webkit-transition:transform .4s cubic-bezier(0.4,0,0.2,1);transition:transform .4s cubic-bezier(0.4,0,0.2,1);-webkit-transition:transform .4s cubic-bezier(0.4,0,0.2,1),-webkit-transform .4s cubic-bezier(0.4,0,0.2,1);transition:transform .4s cubic-bezier(0.4,0,0.2,1),-webkit-transform .4s cubic-bezier(0.4,0,0.2,1);-webkit-box-align:center;box-align:center;-webkit-align-items:center;align-items:center;display:-webkit-box;display:-webkit-flex;display:flex;-webkit-box-orient:vertical;box-orient:vertical;-webkit-flex-direction:column;flex-direction:column;bottom:0;left:0;padding:0 5%;position:absolute;right:0;top:0}.x3wWge,.ONJhl{display:block;height:3em}.eEPege>.x3wWge,.eEPege>.ONJhl{-webkit-box-flex:1;box-flex:1;-webkit-flex-grow:1;flex-grow:1}.J9Nfi{-webkit-flex-shrink:1;flex-shrink:1;max-height:100%}*,*:before,*:after{box-sizing:inherit}html{box-sizing:border-box;-webkit-tap-highlight-color:transparent}body,input,textarea,select,button{color:rgb(32,33,36);font-family:arial,sans-serif}body{background:#fff;direction:ltr;display:-webkit-box;display:-webkit-flex;display:flex;-webkit-box-orient:vertical;-webkit-box-direction:normal;-webkit-flex-direction:column;flex-direction:column;font-size:14px;line-height:1.4286;margin:0;min-height:100vh;padding:0;position:relative}@media (min-width:601px){body{-webkit-box-pack:center;-webkit-justify-content:center;justify-content:center}}[data-style=heading]{color:rgb(32,33,36);font-size:16px;font-weight:500;letter-spacing:.1px;line-height:1.4286}.BDEI9 h2:not(.TrZEUc){color:rgb(32,33,36);font-size:16px;font-weight:500;letter-spacing:.1px;line-height:1.4286}.BDEI9 .fegW5d a:not(.TrZEUc),.BDEI9 .fegW5d button:not(.TrZEUc){color:rgb(25,103,210)}.BDEI9 a{text-decoration:none}.BDEI9 a:not(.TrZEUc),.BDEI9 button:not(.TrZEUc){border-radius:4px;color:rgb(26,115,232);display:inline-block;font-weight:500;letter-spacing:.25px;outline:0;position:relative;z-index:1}.BDEI9 button:not(.TrZEUc){background-color:transparent;cursor:pointer;padding:0;text-align:left}.BDEI9 button:not(.TrZEUc){border:0}.BDEI9 button::-moz-focus-inner{border:0}.BDEI9 a:not(.TrZEUc):focus-visible,.BDEI9 button:not(.TrZEUc):focus-visible{outline:none;position:relative}.BDEI9 a:not(.TrZEUc):focus-visible::after,.BDEI9 button:not(.TrZEUc):focus-visible::after{border:2px solid rgb(24,90,188);border-radius:6px;bottom:-4px;box-shadow:0 0 0 2px rgb(232,240,254);content:"";left:-4px;position:absolute;right:-4px;top:-4px}.BDEI9 a:not(.TrZEUc):focus::after,.BDEI9 a:not(.TrZEUc):active::after,.BDEI9 button:not(.TrZEUc):focus::after,.BDEI9 button:not(.TrZEUc):active::after{background-color:rgba(26,115,232,.15);content:"";position:absolute;z-index:-1}.BDEI9 img:not(.TrZEUc){border:0;max-height:1.3em;vertical-align:middle}@media (min-width:601px){.BDEI9{display:-webkit-box;display:-webkit-flex;display:flex;-webkit-box-orient:vertical;-webkit-box-direction:normal;-webkit-flex-direction:column;flex-direction:column;min-height:100vh;position:relative}.BDEI9::before,.BDEI9::after{-webkit-box-flex:1;-webkit-flex-grow:1;flex-grow:1;content:"";height:24px}.BDEI9::before{min-height:30px}.BDEI9::after{min-height:24px}.BDEI9.LZgQXe::after{min-height:63.9996px}}.gEc4r{display:-webkit-box;display:-webkit-flex;display:flex;height:24px;-webkit-box-pack:center;-webkit-justify-content:center;justify-content:center}.gEc4r.jlqJKb{height:auto;min-height:24px;padding-top:24px}.BivnM{-webkit-box-align:center;-webkit-align-items:center;align-items:center;border-bottom:1px solid #ccc;display:-webkit-box;display:-webkit-flex;display:flex;height:36px;left:0;padding:0 16px;position:absolute;right:0;top:0}.BivnM .ji6sFc{height:14px;margin-right:12px}.O3jdWc{color:rgb(95,99,104);font-size:14px;height:14px;margin-top:-2px}.Zwk8S{display:block;height:37px;width:37px}.wFNE4e{color:rgb(26,115,232)}.HUYFt{display:-webkit-box;display:-webkit-flex;display:flex;-webkit-flex-wrap:wrap;flex-wrap:wrap;font-size:12px;-webkit-box-pack:justify;-webkit-justify-content:space-between;justify-content:space-between;padding:0 24px 14px}@media (min-width:601px){.HUYFt{padding-left:0;padding-right:0;position:absolute;width:100%}}.hXs2T .pUP0Nd{color:rgb(60,64,67)}.hXs2T{margin-left:-16px;margin-right:16px}.N158t{-webkit-appearance:none;appearance:none;background-color:transparent;background-image:url("data:image/svg+xml;base64,PHN2ZyB4bWxucz0iaHR0cDovL3d3dy53My5vcmcvMjAwMC9zdmciIGhlaWdodD0iMjRweCIgdmlld0JveD0iMCAwIDI0IDI0IiB3aWR0aD0iMjRweCIgZmlsbD0iIzQ1NUE2NCI+PHBhdGggZD0iTTAgMGgyNHYyNEgwVjB6IiBmaWxsPSJub25lIi8+PHBhdGggZD0iTTcgMTBsNSA1IDUtNUg3eiIvPjwvc3ZnPg==");background-position:right;background-repeat:no-repeat;border:none;border-radius:4px;color:rgb(95,99,104);cursor:pointer;font-size:12px;line-height:15.9996px;outline:none;padding:16.0002px 24px 16.0002px 16px}.N158t:focus{background-color:rgb(232,234,237)}.M2nKge{list-style:none;margin:0 -16px;padding:0}.vomtoe{display:inline-block;margin:0}.pUP0Nd{background-color:transparent;border-radius:4px;color:rgb(95,99,104);display:inline-block;line-height:15.9996px;outline:none;padding:16px}.pUP0Nd:focus{background-color:rgb(232,234,237)}.pUP0Nd:focus-visible{outline:none;position:relative}.pUP0Nd:focus-visible::after{border:2px solid rgb(24,90,188);border-radius:4px;bottom:-2px;box-shadow:0 0 0 2px rgb(232,240,254);content:"";left:-2px;position:absolute;right:-2px;top:-2px}.JYXaTc{display:-webkit-box;display:-webkit-flex;display:flex;-webkit-box-orient:vertical;-webkit-box-direction:normal;-webkit-flex-direction:column;flex-direction:column;-webkit-box-flex:1;-webkit-flex-grow:1;flex-grow:1;-webkit-flex-wrap:wrap;flex-wrap:wrap;-webkit-box-pack:end;-webkit-justify-content:flex-end;justify-content:flex-end;margin-bottom:-6px;margin-left:-16px;margin-top:32px}.wsArZ[data-ss-mode="1"] .JYXaTc{width:100%}@media (min-width:600px) and (orientation:landscape),all and (min-width:1600px){.NQ5OL .JYXaTc{width:100%}}.JYXaTc.fXx9Lc{margin:0;min-height:0;padding:0}.S1zJGd{-webkit-align-self:flex-start;align-self:flex-start;-webkit-flex-shrink:0;flex-shrink:0;margin-bottom:24px}.O1Slxf{display:-webkit-box;display:-webkit-flex;display:flex;-webkit-box-orient:vertical;-webkit-box-direction:normal;-webkit-flex-direction:row-reverse;flex-direction:row-reverse;-webkit-flex-wrap:wrap;flex-wrap:wrap;width:100%}.TNTaPb,.FO2vFd{display:-webkit-box;display:-webkit-flex;display:flex;-webkit-box-flex:1;-webkit-flex-grow:1;flex-grow:1}@media (min-width:840px){.wsArZ[data-ss-mode="1"] .TNTaPb,.wsArZ[data-ss-mode="1"] .FO2vFd{-webkit-box-flex:unset;-webkit-flex-grow:unset;flex-grow:unset}}@media (min-width:600px) and (orientation:landscape),all and (min-width:1600px){.NQ5OL .JYXaTc:not(.NNItQ) .TNTaPb,.NQ5OL .JYXaTc:not(.NNItQ) .FO2vFd{-webkit-box-flex:unset;-webkit-flex-grow:unset;flex-grow:unset}}.FO2vFd{-webkit-box-pack:flex-start;-webkit-justify-content:flex-start;justify-content:flex-start}.wsArZ[data-ss-mode="1"] .FO2vFd{margin-left:0;margin-right:-16px}@media (min-width:600px) and (orientation:landscape),all and (min-width:1600px){.NQ5OL .FO2vFd{margin-left:0;margin-right:-16px}}.TNTaPb{-webkit-box-pack:flex-end;-webkit-justify-content:flex-end;justify-content:flex-end}.wsArZ[data-ss-mode="1"] .TNTaPb{margin-left:40px;margin-right:0}@media (min-width:600px) and (orientation:landscape),all and (min-width:1600px){.NQ5OL .TNTaPb{margin-left:40px;margin-right:0}}.wsArZ[data-ss-mode="1"] .TNTaPb:empty{margin-left:0;margin-right:0}@media (min-width:600px) and (orientation:landscape),all and (min-width:1600px){.NQ5OL .TNTaPb:empty{margin-left:0;margin-right:0}}.JYXaTc.NNItQ .TNTaPb,.JYXaTc.NNItQ .FO2vFd{-webkit-box-pack:center;-webkit-justify-content:center;justify-content:center}.JYXaTc.NNItQ .TNTaPb,.JYXaTc.F8PBrb .TNTaPb{padding-left:16px}.JYXaTc.F8PBrb .TNTaPb{display:-webkit-box;display:-webkit-flex;display:flex;-webkit-box-pack:justify;-webkit-justify-content:space-between;justify-content:space-between;-webkit-flex-shrink:0;flex-shrink:0;-webkit-flex-wrap:wrap;flex-wrap:wrap;width:100%}.JYXaTc.NNItQ .FO2vFd,.JYXaTc.F8PBrb .TNTaPb+.FO2vFd{margin-top:16px}.JYXaTc:not(.NNItQ) .FO2vFd .mWv92d,.JYXaTc:not(.NNItQ) .FO2vFd .JLt0ke,.JYXaTc:not(.NNItQ) .FO2vFd .J7pUA{text-align:left}.BbN10e{display:block;width:calc(100% - 2px)}.JYXaTc.F8PBrb .O1Slxf{margin:0 -6px;width:calc(100% + 12px)}.JYXaTc.F8PBrb .FO2vFd{margin:0 6px}.o3Yfjb{-webkit-box-flex:1;-webkit-flex-grow:1;flex-grow:1;margin:0 6px;min-width:calc(50% - 12px)}.BbN10e{white-space:nowrap;width:100%}.BbN10e .pIzcPc,.BbN10e .Jskylb{display:block}.mWv92d+.n3Clv,.JLt0ke+.n3Clv{margin-top:32px}.n3Clv .q6oraf{border-radius:16px}.JYXaTc .J7pUA.u3bW4e{background-color:transparent}.J7pUA .snByac{color:#0b57d0;color:var(--gm3-sys-color-primary,#0b57d0);line-height:1.4285714286;margin:16px;text-transform:none}.JYXaTc.JYXaTc .KMdFve{--mdc-ripple-color:var(--gm3-sys-color-on-surface,#1f1f1f);background-color:var(--gm3-sys-color-surface-container,#f0f4f9)}.JYXaTc.JYXaTc .KMdFve .VfPpkd-xl07Ob-ibnC6b-OWXEXe-gk6SMd{background-color:var(--gm3-sys-color-secondary-container,#c2e7ff)}.gNVsKb{color:#1f1f1f;color:var(--gm3-sys-color-on-surface,#1f1f1f)}.J7pUA [jsslot]{margin:0}.BbN10e .pIzcPc,.BbN10e .Jskylb{width:100%}.wsArZ[data-ss-mode="1"] .COi2Ke.lUWEgd.F8PBrb{margin-left:0}@media (min-width:600px) and (orientation:landscape),all and (min-width:1600px){.NQ5OL .COi2Ke.lUWEgd.F8PBrb{margin-left:0}}.wsArZ[data-ss-mode="1"] .COi2Ke.lUWEgd.F8PBrb .TNTaPb{margin-left:0;padding-left:0;width:calc(50% - 24px + 12px)}@media (min-width:600px) and (orientation:landscape),all and (min-width:1600px){.NQ5OL .COi2Ke.lUWEgd.F8PBrb .TNTaPb{margin-left:0;padding-left:0;width:calc(50% - 24px + 12px)}}@media (min-width:840px){.wsArZ[data-ss-mode="1"] .COi2Ke.lUWEgd.F8PBrb .TNTaPb{width:calc(50% - 38px + 12px)}}.COi2Ke.lUWEgd.F8PBrb .FO2vFd{margin-top:2px}.COi2Ke.lUWEgd.F8PBrb .O1Slxf{margin:0 -6px;width:calc(100% + 12px)}.wsArZ[data-ss-mode="1"] .COi2Ke.lUWEgd.F8PBrb .O1Slxf{-webkit-align-self:flex-end;align-self:flex-end;width:100%}@media (min-width:600px) and (orientation:landscape),all and (min-width:1600px){.NQ5OL .COi2Ke.lUWEgd.F8PBrb .O1Slxf{-webkit-align-self:flex-end;align-self:flex-end;width:100%}}.JYXaTc.F8PBrb.lUWEgd.hhh8Yc .FO2vFd{margin-left:10px;margin-right:2px}.wsArZ[data-ss-mode="1"] .JYXaTc.F8PBrb.lUWEgd.hhh8Yc .O1Slxf{-webkit-box-align:end;-webkit-align-items:flex-end;align-items:flex-end;-webkit-box-orient:vertical;-webkit-box-direction:normal;-webkit-flex-flow:column;flex-flow:column}@media (min-width:600px) and (orientation:landscape),all and (min-width:1600px){.NQ5OL .JYXaTc.F8PBrb.lUWEgd.hhh8Yc .O1Slxf{-webkit-box-align:end;-webkit-align-items:flex-end;align-items:flex-end;-webkit-box-orient:vertical;-webkit-box-direction:normal;-webkit-flex-flow:column;flex-flow:column}}.wsArZ[data-ss-mode="1"] .JYXaTc.F8PBrb.lUWEgd.c0e3be .TNTaPb,.wsArZ[data-ss-mode="1"] .JYXaTc.F8PBrb.lUWEgd.c0e3be .FO2vFd{-webkit-box-flex:unset;-webkit-flex-grow:unset;flex-grow:unset}@media (min-width:600px) and (orientation:landscape),all and (min-width:1600px){.NQ5OL .JYXaTc.F8PBrb.lUWEgd.c0e3be .TNTaPb,.NQ5OL .JYXaTc.F8PBrb.lUWEgd.c0e3be .FO2vFd{-webkit-box-flex:unset;-webkit-flex-grow:unset;flex-grow:unset}}.JYXaTc.F8PBrb.lUWEgd.c0e3be.NNItQ .TNTaPb{width:100%}.JYXaTc.F8PBrb.lUWEgd.c0e3be .FO2vFd{-webkit-box-pack:center;-webkit-justify-content:center;justify-content:center;padding-left:16px}.wsArZ[data-ss-mode="1"] .JYXaTc.F8PBrb.lUWEgd.c0e3be .FO2vFd{-webkit-box-pack:start;-webkit-justify-content:flex-start;justify-content:flex-start;margin-top:0;margin-right:6px;padding-left:0}@media (min-width:600px) and (orientation:landscape),all and (min-width:1600px){.NQ5OL .JYXaTc.F8PBrb.lUWEgd.c0e3be .FO2vFd{-webkit-box-pack:start;-webkit-justify-content:flex-start;justify-content:flex-start;margin-top:0;margin-right:6px;padding-left:0}}.JYXaTc.F8PBrb.lUWEgd.c0e3be.NNItQ .O1Slxf{-webkit-box-align:center;-webkit-align-items:center;align-items:center;-webkit-box-orient:vertical;-webkit-box-direction:normal;-webkit-flex-flow:column;flex-flow:column}.wsArZ[data-ss-mode="1"] .JYXaTc.F8PBrb.lUWEgd.c0e3be.NNItQ .O1Slxf{width:calc(50% - 24px + 12px)}@media (min-width:600px) and (orientation:landscape),all and (min-width:1600px){.NQ5OL .JYXaTc.F8PBrb.lUWEgd.c0e3be.NNItQ .O1Slxf{width:calc(50% - 24px + 12px)}}@media (min-width:840px){.wsArZ[data-ss-mode="1"] .JYXaTc.F8PBrb.lUWEgd.c0e3be.NNItQ .O1Slxf{width:calc(50% - 38px + 12px)}}.JYXaTc.F8PBrb.lUWEgd.x8Ikx .TNTaPb,.JYXaTc.F8PBrb.lUWEgd.N0osAb .TNTaPb{-webkit-box-orient:vertical;-webkit-box-direction:normal;-webkit-flex-flow:column;flex-flow:column}.wsArZ[data-ss-mode="1"] .JYXaTc.F8PBrb.lUWEgd.x8Ikx .TNTaPb,.wsArZ[data-ss-mode="1"] .JYXaTc.F8PBrb.lUWEgd.N0osAb .TNTaPb{width:100%}@media (min-width:600px) and (orientation:landscape),all and (min-width:1600px){.NQ5OL .JYXaTc.F8PBrb.lUWEgd.x8Ikx .TNTaPb,.NQ5OL .JYXaTc.F8PBrb.lUWEgd.N0osAb .TNTaPb{width:100%}}.JYXaTc.F8PBrb.lUWEgd.x8Ikx .FO2vFd,.JYXaTc.F8PBrb.lUWEgd.N0osAb .FO2vFd{-webkit-box-pack:center;-webkit-justify-content:center;justify-content:center;margin-left:16px;margin-right:2px;margin-top:0}.wsArZ[data-ss-mode="1"] .JYXaTc.F8PBrb.lUWEgd.x8Ikx .FO2vFd,.wsArZ[data-ss-mode="1"] .JYXaTc.F8PBrb.lUWEgd.N0osAb .FO2vFd{margin-left:0}@media (min-width:600px) and (orientation:landscape),all and (min-width:1600px){.NQ5OL .JYXaTc.F8PBrb.lUWEgd.x8Ikx .FO2vFd,.NQ5OL .JYXaTc.F8PBrb.lUWEgd.N0osAb .FO2vFd{margin-left:0}}.JYXaTc.F8PBrb.lUWEgd.x8Ikx .O1Slxf,.JYXaTc.F8PBrb.lUWEgd.N0osAb .O1Slxf{-webkit-box-align:center;-webkit-align-items:center;align-items:center;-webkit-box-orient:vertical;-webkit-box-direction:normal;-webkit-flex-flow:column;flex-flow:column}.wsArZ[data-ss-mode="1"] .JYXaTc.F8PBrb.lUWEgd.x8Ikx .O1Slxf,.wsArZ[data-ss-mode="1"] .JYXaTc.F8PBrb.lUWEgd.N0osAb .O1Slxf{width:calc(50% - 24px + 12px)}@media (min-width:600px) and (orientation:landscape),all and (min-width:1600px){.NQ5OL .JYXaTc.F8PBrb.lUWEgd.x8Ikx .O1Slxf,.NQ5OL .JYXaTc.F8PBrb.lUWEgd.N0osAb .O1Slxf{width:calc(50% - 24px + 12px)}}@media (min-width:840px){.wsArZ[data-ss-mode="1"] .JYXaTc.F8PBrb.lUWEgd.x8Ikx .O1Slxf,.wsArZ[data-ss-mode="1"] .JYXaTc.F8PBrb.lUWEgd.N0osAb .O1Slxf{width:calc(50% - 38px + 12px)}}.JYXaTc.F8PBrb.lUWEgd.N0osAb .FO2vFd{margin:0;padding-left:16px;width:calc(100% - 12px)}.wsArZ[data-ss-mode="1"] .JYXaTc.F8PBrb.lUWEgd.N0osAb .FO2vFd{padding-left:0}@media (min-width:600px) and (orientation:landscape),all and (min-width:1600px){.NQ5OL .JYXaTc.F8PBrb.lUWEgd.N0osAb .FO2vFd{padding-left:0}}.JYXaTc.F8PBrb.N0osAb .mWv92d,.JYXaTc.F8PBrb.N0osAb .mWv92d .pIzcPc{display:block;width:100%}.JYXaTc.F8PBrb.lUWEgd.N0osAb .BbN10e .Jskylb,.JYXaTc.F8PBrb.lUWEgd.N0osAb .mWv92d .pIzcPc{margin-top:4px;margin-bottom:4px}.wsArZ[data-ss-mode="1"] .JYXaTc.F8PBrb{margin-left:0}@media (min-width:600px) and (orientation:landscape),all and (min-width:1600px){.NQ5OL .JYXaTc.F8PBrb{margin-left:0}}.wsArZ[data-ss-mode="1"] .JYXaTc.F8PBrb .TNTaPb{-webkit-box-flex:unset;-webkit-flex-grow:unset;flex-grow:unset;margin-left:0;padding-left:0;width:calc(50% - 24px + 12px)}@media (min-width:600px) and (orientation:landscape),all and (min-width:1600px){.NQ5OL .JYXaTc.F8PBrb .TNTaPb{-webkit-box-flex:unset;-webkit-flex-grow:unset;flex-grow:unset;margin-left:0;padding-left:0;width:calc(50% - 24px + 12px)}}@media (min-width:840px){.wsArZ[data-ss-mode="1"] .JYXaTc.F8PBrb .TNTaPb{width:calc(50% - 38px + 12px)}}.JYXaTc.F8PBrb.NNItQ .TNTaPb{width:100%}.JYXaTc.F8PBrb .FO2vFd{margin-left:6px;margin-right:6px}.wsArZ[data-ss-mode="1"] .JYXaTc.F8PBrb .FO2vFd{margin-left:2px}@media (min-width:600px) and (orientation:landscape),all and (min-width:1600px){.NQ5OL .JYXaTc.F8PBrb .FO2vFd{margin-left:2px}}.JYXaTc.F8PBrb .O1Slxf{-webkit-box-align:start;-webkit-align-items:flex-start;align-items:flex-start;-webkit-box-orient:vertical;-webkit-box-direction:normal;-webkit-flex-direction:column;flex-direction:column;margin:0 -6px;width:calc(100% + 12px)}.wsArZ[data-ss-mode="1"] .JYXaTc.F8PBrb .O1Slxf{-webkit-box-align:end;-webkit-align-items:flex-end;align-items:flex-end;-webkit-align-self:flex-end;align-self:flex-end;width:100%}@media (min-width:600px) and (orientation:landscape),all and (min-width:1600px){.NQ5OL .JYXaTc.F8PBrb .O1Slxf{-webkit-box-align:end;-webkit-align-items:flex-end;align-items:flex-end;-webkit-align-self:flex-end;align-self:flex-end;width:100%}}.JYXaTc.F8PBrb.NNItQ .O1Slxf{-webkit-box-align:center;-webkit-align-items:center;align-items:center}.wsArZ[data-ss-mode="1"] .JYXaTc.F8PBrb.NNItQ .O1Slxf{width:calc(50% - 24px + 12px)}@media (min-width:600px) and (orientation:landscape),all and (min-width:1600px){.NQ5OL .JYXaTc.F8PBrb.NNItQ .O1Slxf{width:calc(50% - 24px + 12px)}}@media (min-width:840px){.wsArZ[data-ss-mode="1"] .JYXaTc.F8PBrb.NNItQ .O1Slxf{width:calc(50% - 38px + 12px)}}.COi2Ke.lUWEgd.F8PBrb .FO2vFd{margin-right:2px}.JYXaTc.F8PBrb.lUWEgd.c0e3be .FO2vFd{margin-left:2px}.JYXaTc.F8PBrb.lUWEgd.c0e3be .O1Slxf{-webkit-box-orient:horizontal;-webkit-box-direction:reverse;-webkit-flex-direction:row-reverse;flex-direction:row-reverse}.ObDc3{display:-webkit-box;display:-webkit-flex;display:flex;-webkit-box-orient:vertical;-webkit-box-direction:normal;-webkit-flex-direction:column;flex-direction:column;margin-bottom:32px}@media (min-width:840px){.ObDc3{margin-bottom:32px}}.wsArZ[data-ss-mode="1"] .ObDc3{margin-bottom:0}@media (min-width:600px) and (orientation:landscape),all and (min-width:1600px){.NQ5OL .ObDc3{margin-bottom:0}}.Su9bff{-webkit-box-align:center;-webkit-align-items:center;align-items:center;text-align:center}.vAV9bf{color:#1f1f1f;color:var(--gm3-sys-color-on-surface,#1f1f1f);font-family:"Google Sans",roboto,"Noto Sans Myanmar UI",arial,sans-serif;font-weight:400;font-weight:var(--c-tfwt,400);line-height:1.25;margin-bottom:0;margin-bottom:var(--c-ts-b,0);margin-top:24px;margin-top:var(--c-ts-t,24px);word-break:break-word;font-size:2rem;font-size:var(--wf-tfs,2rem)}@media (min-width:840px){.vAV9bf{line-height:1.2222222222;font-size:2.25rem;font-size:var(--wf-tfs-bp3,2.25rem)}}@media (min-width:960px){.vAV9bf{line-height:1.2222222222;font-size:2.25rem;font-size:var(--wf-tfs-bp3,2.25rem)}}@media (min-width:1600px){.vAV9bf{line-height:1.1818181818;font-size:2.75rem;font-size:var(--wf-tfs-bp5,2.75rem)}}.gNJDp{color:#1f1f1f;color:var(--gm3-sys-color-on-surface,#1f1f1f);font-family:"Google Sans",roboto,"Noto Sans Myanmar UI",arial,sans-serif;font-weight:400;font-weight:var(--c-stfwt,400);letter-spacing:0rem;line-height:1.5;margin-bottom:0;margin-bottom:var(--c-sts-b,0);margin-top:16px;margin-top:var(--c-sts-t,16px);font-size:1rem;font-size:var(--wf-stfs,1rem)}@media (min-width:1600px){.gNJDp{line-height:1.5;font-size:1rem;font-size:var(--wf-stfs-bp5,1rem)}}.gNJDp:empty{display:none}.I7GnLc{font-weight:500;letter-spacing:.25px;min-height:24px}.SOeSgb{height:32px}.I7GnLc,.SOeSgb{margin-bottom:0;margin-bottom:var(--c-sts-b,0);margin-top:16px;margin-top:var(--c-sts-t,16px)}.ObDc3.ZYOIke .I7GnLc,.ObDc3.ZYOIke .SOeSgb{margin-bottom:0;margin-top:16px}.SfkAJe{-webkit-box-flex:1;-webkit-flex-grow:1;flex-grow:1}.sQecwc{display:hidden}*,*::before,*::after{box-sizing:inherit}html{box-sizing:border-box;-webkit-tap-highlight-color:rgba(0,0,0,0)}.jR8x9d{color-scheme:light}.jR8x9d,.jR8x9d input,.jR8x9d textarea,.jR8x9d select,.jR8x9d button{color:#1f1f1f;color:var(--gm3-sys-color-on-surface,#1f1f1f);font-family:"Google Sans",roboto,"Noto Sans Myanmar UI",arial,sans-serif}.jR8x9d{background-color:#fff;background-color:var(--gm3-sys-color-surface-container-lowest,#fff);direction:ltr;font-size:0.875rem;font-weight:400;letter-spacing:0rem;line-height:1.4285714286;margin:0;padding:0}.jR8x9d [data-style=heading]{color:#1f1f1f;color:var(--gm3-sys-color-on-surface,#1f1f1f);font-family:"Google Sans",roboto,"Noto Sans Myanmar UI",arial,sans-serif;font-size:1.25rem;font-weight:400;letter-spacing:0rem;line-height:1.2}.S7xv8{display:-webkit-box;display:-webkit-flex;display:flex;-webkit-box-orient:vertical;-webkit-box-direction:normal;-webkit-flex-direction:column;flex-direction:column;min-height:100vh;background:#fff;background:var(--gm3-sys-color-surface-container-lowest,#fff);-webkit-box-pack:justify;-webkit-justify-content:space-between;justify-content:space-between;padding:0}@media (min-width:600px){.S7xv8{background:#f0f4f9;background:var(--gm3-sys-color-surface-container,#f0f4f9);-webkit-box-pack:center;-webkit-justify-content:center;justify-content:center;padding:48px 0}}@media (min-width:600px) and (orientation:landscape){.S7xv8{background:#fff;background:var(--gm3-sys-color-surface-container-lowest,#fff);-webkit-box-pack:justify;-webkit-justify-content:space-between;justify-content:space-between;padding:0}}@media (min-width:960px) and (orientation:landscape){.S7xv8{background:#f0f4f9;background:var(--gm3-sys-color-surface-container,#f0f4f9);-webkit-box-pack:center;-webkit-justify-content:center;justify-content:center;padding:48px 0}}.fAlnEc a:not(.TrZEUc):not(.WpHeLc){outline-offset:2px;text-decoration:none}.fAlnEc a:not(.TrZEUc):not(.WpHeLc):hover{text-decoration:underline}.fAlnEc button:not(.TrZEUc){background-color:transparent;border:0;cursor:pointer;font-size:inherit;outline:none;padding:0;position:relative;text-align:left}.fAlnEc a:not(.TrZEUc):not(.WpHeLc),.fAlnEc button:not(.TrZEUc){color:#0b57d0;color:var(--gm3-sys-color-primary,#0b57d0);border-radius:4px;font-weight:500;letter-spacing:0.015625rem;z-index:1}.fAlnEc a:not(.TrZEUc):not(.WpHeLc):focus-visible{outline:2px solid #0b57d0;outline:2px solid var(--gm3-sys-color-primary,#0b57d0)}.fAlnEc .gNJDp a:not(.TrZEUc):not(.WpHeLc),.fAlnEc .gNJDp button:not(.TrZEUc){font-weight:500;font-weight:var(--c-stfwt,500)}.fAlnEc .PsAlOe a:not(.TrZEUc),.fAlnEc .PsAlOe button:not(.TrZEUc){text-decoration:underline}.fAlnEc .PsAlOe.sj692e a:not(.TrZEUc),.fAlnEc .PsAlOe.sj692e button:not(.TrZEUc){color:#0842a0;color:var(--gm3-sys-color-on-primary-container,#0842a0)}.fAlnEc .Su9bff a:not(.L3JCSb),.fAlnEc .Su9bff button:not(.L3JCSb){text-align:center}.fAlnEc .PsAlOe.Xq8bDe a:not(.TrZEUc),.fAlnEc .PsAlOe.Xq8bDe button:not(.TrZEUc){color:#410e0b;color:var(--gm3-sys-color-on-error-container,#8c1d18)}.fAlnEc .PsAlOe.rNe0id a:not(.TrZEUc),.fAlnEc .PsAlOe.rNe0id button:not(.TrZEUc){color:var(--wf-color-warning-text,#421f00)}.fAlnEc .PsAlOe.YFdWic a:not(.TrZEUc),.fAlnEc .PsAlOe.YFdWic button:not(.TrZEUc){color:#444746;color:var(--gm3-sys-color-on-surface-variant,#444746)}.fAlnEc button:not(.TrZEUc)::-moz-focus-inner{border:0}.fAlnEc button:not(.TrZEUc):focus-visible::after{border:2px solid;border-color:#0b57d0;border-color:var(--gm3-sys-color-primary,#0b57d0);box-shadow:0 0 0 2px #d3e3fd;box-shadow:0 0 0 2px var(--gm3-sys-color-primary-container,#d3e3fd);border-radius:12px;content:"";position:absolute;pointer-events:none;inset:-9px;bottom:-5px;top:-5px}.fAlnEc button:not(.TrZEUc)::before{background-color:#0b57d0;background-color:var(--gm3-sys-color-primary,#0b57d0);border-radius:8px;bottom:-1px;content:"";left:-5px;opacity:0;pointer-events:none;position:absolute;right:-5px;top:-1px;z-index:-1}.fAlnEc button:not(.TrZEUc):hover::before{opacity:.08}.fAlnEc button:not(.TrZEUc):focus::before,.fAlnEc button:not(.TrZEUc):active::before{opacity:.1}.fAlnEc img:not(.TrZEUc){border:0;max-height:1.3em;vertical-align:middle}@media screen and (prefers-color-scheme:dark){.jR8x9d{color-scheme:dark}.jR8x9d .Y5O54e{display:-webkit-inline-box;display:-webkit-inline-flex;display:inline-flex;position:relative}.jR8x9d .Y5O54e[hidden]{display:none}.jR8x9d .Y5O54e .UMrnmb-lP5Lpb-yrriRe{width:inherit}.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b{padding-left:16px;padding-right:16px}[dir=rtl] .jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b,.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b[dir=rtl]{padding-left:16px;padding-right:16px}.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-f7MjDc{margin-left:0;margin-right:8px}[dir=rtl] .jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-f7MjDc,.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-f7MjDc[dir=rtl]{margin-left:8px;margin-right:0}.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb.UMrnmb-h0T7hb-M1Soyc-Bz112c .VfPpkd-StrnGf-rymPhb-ibnC6b{padding-left:48px;padding-right:16px}[dir=rtl] .jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb.UMrnmb-h0T7hb-M1Soyc-Bz112c .VfPpkd-StrnGf-rymPhb-ibnC6b,.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb.UMrnmb-h0T7hb-M1Soyc-Bz112c .VfPpkd-StrnGf-rymPhb-ibnC6b[dir=rtl]{padding-left:16px;padding-right:48px}.jR8x9d .Y5O54e .VfPpkd-xl07Ob-XxIAqe-OWXEXe-uxVfW-FNFY6c-uFfGwd{border-top-left-radius:0;border-top-right-radius:0}.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe:hover .VfPpkd-fmcmS-OyKIhb::before,.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-fmcmS-OyKIhb::before{opacity:.08;opacity:var(--mdc-ripple-hover-opacity,.08)}.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-fmcmS-OyKIhb::before,.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-fmcmS-OyKIhb::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:0;opacity:var(--mdc-ripple-focus-opacity,0)}.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe .VfPpkd-fmcmS-OyKIhb::before,.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe .VfPpkd-fmcmS-OyKIhb::after{background-color:rgb(241,243,244);background-color:var(--mdc-ripple-color,rgb(241,243,244))}.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd,.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me)+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd{color:rgb(154,160,166)}.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe .VfPpkd-fmcmS-wGMbrd{caret-color:rgb(138,180,248)}.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-wGMbrd{color:rgb(232,234,237)}.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me){background-color:rgb(60,64,67)}.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me)+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-W0vJo-fmcmS{color:rgb(154,160,166)}.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(189,193,198)}.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe:hover:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(248,249,250)}.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe:hover:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgb(248,249,250)}.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgb(154,160,166)}.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::after{border-bottom-color:rgb(138,180,248)}}@media screen and (prefers-color-scheme:dark){.boqAccountsWireframeThemesMaterialnextBaseBodyEl .GmFilledAutocompleteDarkTheme .mdc-text-field:not(.mdc-text-field--disabled) .mdc-text-field__input::-webkit-input-placeholder{color:rgb(189,193,198)}.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-wGMbrd::placeholder{color:rgb(189,193,198)}}@media screen and (prefers-color-scheme:dark){.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-wGMbrd:-ms-input-placeholder{color:rgb(189,193,198)}.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-MvKemf-OWXEXe-qdIk2c{color:rgb(154,160,166)}.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-MvKemf-OWXEXe-iJ4yB{color:rgb(154,160,166)}.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc{color:rgb(154,160,166)}.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-UbuQg{color:rgb(154,160,166)}.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-wGMbrd{color:rgba(232,234,237,.38)}.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me{background-color:rgba(232,234,237,.04)}.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgba(232,234,237,.38)}.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-NLUYnc-V67aGc,.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc,.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-TvZj5c-OWXEXe-UbuQg,.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-W0vJo-fmcmS,.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd,.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd{color:rgba(232,234,237,.38)}}@media screen and (prefers-color-scheme:dark){.boqAccountsWireframeThemesMaterialnextBaseBodyEl .GmFilledAutocompleteDarkTheme .mdc-text-field.mdc-text-field--disabled .mdc-text-field__input::-webkit-input-placeholder{color:rgba(232,234,237,.38)}.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-wGMbrd::placeholder{color:rgba(232,234,237,.38)}}@media screen and (prefers-color-scheme:dark){.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-wGMbrd:-ms-input-placeholder{color:rgba(232,234,237,.38)}.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-MvKemf-OWXEXe-qdIk2c,.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-MvKemf-OWXEXe-iJ4yB{color:rgba(232,234,237,.38)}.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(138,180,248)}.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc .VfPpkd-fmcmS-wGMbrd{caret-color:rgb(246,174,169)}.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me)+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-W0vJo-fmcmS{color:rgb(242,139,130)}.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-UbuQg{color:rgb(242,139,130)}.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgb(246,174,169)}.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::after{border-bottom-color:rgb(246,174,169)}.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:hover:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(246,174,169)}.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:hover:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me)+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-W0vJo-fmcmS{color:rgb(246,174,169)}.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:hover:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-UbuQg{color:rgb(246,174,169)}.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:hover:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgb(246,174,169)}.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc{color:rgb(138,180,248)}.jR8x9d .Y5O54e .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(246,174,169)}.jR8x9d .Y5O54e .VfPpkd-xl07Ob-XxIAqe{box-shadow:0 2px 1px -1px rgba(0,0,0,.2),0 1px 1px 0 rgba(0,0,0,.14),0 1px 3px 0 rgba(0,0,0,.12);background-color:rgb(32,33,36)}.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb{font-family:Roboto,Arial,sans-serif;line-height:1.5rem;font-size:1rem;letter-spacing:.00625em;font-weight:400;color:rgb(232,234,237);position:relative}.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-IhFlZd{color:rgb(154,160,166)}.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS{color:rgb(232,234,237)}.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c{opacity:.38}.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd,.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b,.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-f7MjDc,.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-f7MjDc{color:rgb(232,234,237)}.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:0}.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd{background-color:rgba(138,180,248,.24)}.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before,.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::after{background-color:rgb(138,180,248);background-color:var(--mdc-ripple-color,rgb(138,180,248))}.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before,.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before,.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS{color:rgb(154,160,166)}.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic{border-bottom-color:rgba(232,234,237,.12)}.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc{color:rgb(232,234,237)}.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-pZXsl::before,.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-pZXsl::after{background-color:rgb(232,234,237);background-color:var(--mdc-ripple-color,rgb(232,234,237))}.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before,.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before,.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}}@media screen and (prefers-color-scheme:dark) and (-ms-high-contrast:active),screen and (prefers-color-scheme:dark) and (forced-colors:active){.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS{color:GrayText}.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c{opacity:1}}@media screen and (prefers-color-scheme:dark){.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb .VfPpkd-BFbNVe-bF1uUb{width:100%;height:100%;top:0;left:0}.jR8x9d .Y5O54e .VfPpkd-StrnGf-rymPhb .VfPpkd-BFbNVe-bF1uUb{opacity:.08}.jR8x9d .NGdKgb{display:-webkit-inline-box;display:-webkit-inline-flex;display:inline-flex;position:relative}.jR8x9d .NGdKgb[hidden]{display:none}.jR8x9d .NGdKgb .UMrnmb-lP5Lpb-yrriRe{width:inherit}.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b{padding-left:16px;padding-right:16px}[dir=rtl] .jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b,.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b[dir=rtl]{padding-left:16px;padding-right:16px}.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-f7MjDc{margin-left:0;margin-right:8px}[dir=rtl] .jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-f7MjDc,.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb.VfPpkd-StrnGf-rymPhb-OWXEXe-Bz112c-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-f7MjDc[dir=rtl]{margin-left:8px;margin-right:0}.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb.UMrnmb-h0T7hb-M1Soyc-Bz112c .VfPpkd-StrnGf-rymPhb-ibnC6b{padding-left:48px;padding-right:16px}[dir=rtl] .jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb.UMrnmb-h0T7hb-M1Soyc-Bz112c .VfPpkd-StrnGf-rymPhb-ibnC6b,.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb.UMrnmb-h0T7hb-M1Soyc-Bz112c .VfPpkd-StrnGf-rymPhb-ibnC6b[dir=rtl]{padding-left:16px;padding-right:48px}.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-wGMbrd{color:rgb(232,234,237);color:var(--gm-outlinedtextfield-ink-color,rgb(232,234,237))}.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe .VfPpkd-fmcmS-wGMbrd{caret-color:rgb(138,180,248);caret-color:var(--gm-outlinedtextfield-caret-color,rgb(138,180,248))}.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me)+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-W0vJo-fmcmS{color:rgb(154,160,166);color:var(--gm-outlinedtextfield-helper-text-color,rgb(154,160,166))}.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd,.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me)+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd{color:rgb(154,160,166)}.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(154,160,166);color:var(--gm-outlinedtextfield-label-color,rgb(154,160,166))}.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe:hover:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(248,249,250)}.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Brv4Fb,.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Ra9xwd,.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-MpmGFe{border-color:rgb(189,193,198);border-color:var(--gm-outlinedtextfield-outline-color,rgb(189,193,198))}.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Brv4Fb,.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Ra9xwd,.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-MpmGFe{border-color:rgb(248,249,250)}}@media screen and (prefers-color-scheme:dark){.boqAccountsWireframeThemesMaterialnextBaseBodyEl .GmOutlinedAutocompleteDarkTheme .mdc-text-field:not(.mdc-text-field--disabled) .mdc-text-field__input::-webkit-input-placeholder{color:rgb(189,193,198);color:var(--gm-outlinedtextfield-placeholder-color,rgb(189,193,198))}.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-wGMbrd::placeholder{color:rgb(189,193,198);color:var(--gm-outlinedtextfield-placeholder-color,rgb(189,193,198))}}@media screen and (prefers-color-scheme:dark){.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-wGMbrd:-ms-input-placeholder{color:rgb(189,193,198);color:var(--gm-outlinedtextfield-placeholder-color,rgb(189,193,198))}.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-MvKemf-OWXEXe-qdIk2c{color:rgb(154,160,166);color:var(--gm-outlinedtextfield-prefix-color,rgb(154,160,166))}.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-MvKemf-OWXEXe-iJ4yB{color:rgb(154,160,166);color:var(--gm-outlinedtextfield-suffix-color,rgb(154,160,166))}.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc{color:rgb(154,160,166)}.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-UbuQg{color:rgb(154,160,166)}.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-wGMbrd{color:rgba(232,234,237,.38);color:var(--gm-outlinedtextfield-ink-color--disabled,rgba(232,234,237,.38))}.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-NSFCdd-Brv4Fb,.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-NSFCdd-Ra9xwd,.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-NSFCdd-MpmGFe{border-color:rgba(232,234,237,.12);border-color:var(--gm-outlinedtextfield-outline-color--disabled,rgba(232,234,237,.12))}.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-NLUYnc-V67aGc{color:rgba(232,234,237,.38);color:var(--gm-outlinedtextfield-label-color--disabled,rgba(232,234,237,.38))}.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc{color:rgba(232,234,237,.38);color:var(--gm-outlinedtextfield-icon-color--disabled,rgba(232,234,237,.38))}.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-TvZj5c-OWXEXe-UbuQg{color:rgba(232,234,237,.38);color:var(--gm-outlinedtextfield-icon-color--disabled,rgba(232,234,237,.38))}.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-W0vJo-fmcmS{color:rgba(232,234,237,.38);color:var(--gm-outlinedtextfield-helper-text-color--disabled,rgba(232,234,237,.38))}.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd,.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd{color:rgba(232,234,237,.38);color:var(--gm-outlinedtextfield-character-counter-color--disabled,rgba(232,234,237,.38))}}@media screen and (prefers-color-scheme:dark){.boqAccountsWireframeThemesMaterialnextBaseBodyEl .GmOutlinedAutocompleteDarkTheme .mdc-text-field.mdc-text-field--disabled .mdc-text-field__input::-webkit-input-placeholder{color:rgba(232,234,237,.38);color:var(--gm-outlinedtextfield-placeholder-color--disabled,rgba(232,234,237,.38))}.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-wGMbrd::placeholder{color:rgba(232,234,237,.38);color:var(--gm-outlinedtextfield-placeholder-color--disabled,rgba(232,234,237,.38))}}@media screen and (prefers-color-scheme:dark){.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-wGMbrd:-ms-input-placeholder{color:rgba(232,234,237,.38);color:var(--gm-outlinedtextfield-placeholder-color--disabled,rgba(232,234,237,.38))}.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-MvKemf-OWXEXe-qdIk2c{color:rgba(232,234,237,.38);color:var(--gm-outlinedtextfield-prefix-color--disabled,rgba(232,234,237,.38))}.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-MvKemf-OWXEXe-iJ4yB{color:rgba(232,234,237,.38);color:var(--gm-outlinedtextfield-suffix-color--disabled,rgba(232,234,237,.38))}.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Brv4Fb,.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Ra9xwd,.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-MpmGFe{border-color:rgb(138,180,248);border-color:var(--gm-outlinedtextfield-outline-color--stateful,rgb(138,180,248))}.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(138,180,248);color:var(--gm-outlinedtextfield-label-color--stateful,rgb(138,180,248))}.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc .VfPpkd-fmcmS-wGMbrd{caret-color:rgb(242,139,130);caret-color:var(--gm-outlinedtextfield-caret-color--error,rgb(242,139,130))}.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me)+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-W0vJo-fmcmS{color:rgb(242,139,130);color:var(--gm-outlinedtextfield-helper-text-color--error,rgb(242,139,130))}.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:hover:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me)+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-W0vJo-fmcmS{color:rgb(246,174,169)}.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:hover:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(246,174,169)}.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:hover:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-UbuQg{color:rgb(246,174,169)}.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Brv4Fb,.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Ra9xwd,.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-MpmGFe{border-color:rgb(246,174,169)}.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Brv4Fb,.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Ra9xwd,.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-MpmGFe{border-color:rgb(242,139,130);border-color:var(--gm-outlinedtextfield-outline-color--error,rgb(242,139,130))}.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-UbuQg{color:rgb(242,139,130);color:var(--gm-outlinedtextfield-icon-color--error,rgb(242,139,130))}.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Brv4Fb,.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Ra9xwd,.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-MpmGFe{border-color:rgb(242,139,130);border-color:var(--gm-outlinedtextfield-outline-color--error-stateful,rgb(242,139,130))}.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc{color:rgb(138,180,248);color:var(--gm-outlinedtextfield-label-color--stateful,rgb(138,180,248))}.jR8x9d .NGdKgb .VfPpkd-fmcmS-yrriRe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(242,139,130);color:var(--gm-outlinedtextfield-label-color--error,rgb(242,139,130))}.jR8x9d .NGdKgb .VfPpkd-xl07Ob-XxIAqe{box-shadow:0 2px 1px -1px rgba(0,0,0,.2),0 1px 1px 0 rgba(0,0,0,.14),0 1px 3px 0 rgba(0,0,0,.12);background-color:rgb(32,33,36);margin-bottom:8px}.jR8x9d .NGdKgb.UMrnmb-h0T7hb-OWXEXe-di8rgd-V67aGc .VfPpkd-xl07Ob-XxIAqe,.jR8x9d .NGdKgb .VfPpkd-xl07Ob-XxIAqe-OWXEXe-uxVfW-FNFY6c-uFfGwd{margin-bottom:0}.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb{font-family:Roboto,Arial,sans-serif;line-height:1.5rem;font-size:1rem;letter-spacing:.00625em;font-weight:400;color:rgb(232,234,237);position:relative}.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-IhFlZd{color:rgb(154,160,166)}.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS{color:rgb(232,234,237)}.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c{opacity:.38}.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd,.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b,.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-f7MjDc,.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-f7MjDc{color:rgb(232,234,237)}.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:0}.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd{background-color:rgba(138,180,248,.24)}.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before,.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::after{background-color:rgb(138,180,248);background-color:var(--mdc-ripple-color,rgb(138,180,248))}.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before,.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before,.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS{color:rgb(154,160,166)}.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic{border-bottom-color:rgba(232,234,237,.12)}.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc{color:rgb(232,234,237)}.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-pZXsl::before,.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-pZXsl::after{background-color:rgb(232,234,237);background-color:var(--mdc-ripple-color,rgb(232,234,237))}.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before,.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before,.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}}@media screen and (prefers-color-scheme:dark) and (-ms-high-contrast:active),screen and (prefers-color-scheme:dark) and (forced-colors:active){.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS{color:GrayText}.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c{opacity:1}}@media screen and (prefers-color-scheme:dark){.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb .VfPpkd-BFbNVe-bF1uUb{width:100%;height:100%;top:0;left:0}.jR8x9d .NGdKgb .VfPpkd-StrnGf-rymPhb .VfPpkd-BFbNVe-bF1uUb{opacity:.08}.jR8x9d .DUonjc{background-color:rgb(32,33,36);border-bottom-color:rgb(95,99,104)}.jR8x9d .DUonjc .VfPpkd-WLXbod{background-color:rgb(32,33,36)}.jR8x9d .DUonjc .VfPpkd-Rj7Y9b{color:rgb(232,234,237)}.jR8x9d .DUonjc .VfPpkd-WLXbod{border-bottom-color:rgb(95,99,104)}.jR8x9d .DUonjc .VfPpkd-r7nwK{color:rgb(32,33,36)}.jR8x9d .DUonjc .VfPpkd-r7nwK{background-color:rgb(138,180,248)}.jR8x9d .DUonjc .VfPpkd-LgbsSe:not(:disabled){background-color:transparent}.jR8x9d .DUonjc .VfPpkd-LgbsSe:not(:disabled){color:rgb(138,180,248);color:var(--gm-colortextbutton-ink-color,rgb(138,180,248))}.jR8x9d .DUonjc .VfPpkd-LgbsSe:disabled{color:rgba(232,234,237,.38);color:var(--gm-colortextbutton-disabled-ink-color,rgba(232,234,237,.38))}.jR8x9d .DUonjc .VfPpkd-LgbsSe .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo,.jR8x9d .DUonjc .VfPpkd-LgbsSe .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:rgb(138,180,248)}}@media screen and (prefers-color-scheme:dark) and (-ms-high-contrast:active),screen and (prefers-color-scheme:dark) and (forced-colors:active){.jR8x9d .DUonjc .VfPpkd-LgbsSe .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo,.jR8x9d .DUonjc .VfPpkd-LgbsSe .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:CanvasText}}@media screen and (prefers-color-scheme:dark){.jR8x9d .DUonjc .VfPpkd-LgbsSe:hover:not(:disabled),.jR8x9d .DUonjc .VfPpkd-LgbsSe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:disabled),.jR8x9d .DUonjc .VfPpkd-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d):focus:not(:disabled),.jR8x9d .DUonjc .VfPpkd-LgbsSe:active:not(:disabled){color:rgb(174,203,250);color:var(--gm-colortextbutton-ink-color--stateful,rgb(174,203,250))}.jR8x9d .DUonjc .VfPpkd-LgbsSe .VfPpkd-Jh9lGc::before,.jR8x9d .DUonjc .VfPpkd-LgbsSe .VfPpkd-Jh9lGc::after{background-color:rgb(174,203,250);background-color:var(--gm-colortextbutton-state-color,rgb(174,203,250))}.jR8x9d .DUonjc .VfPpkd-LgbsSe:hover .VfPpkd-Jh9lGc::before,.jR8x9d .DUonjc .VfPpkd-LgbsSe.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.jR8x9d .DUonjc .VfPpkd-LgbsSe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.jR8x9d .DUonjc .VfPpkd-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.jR8x9d .DUonjc .VfPpkd-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .DUonjc .VfPpkd-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.jR8x9d .DUonjc .VfPpkd-LgbsSe.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}.jR8x9d .DUonjc .VfPpkd-LgbsSe:disabled:hover .VfPpkd-Jh9lGc::before,.jR8x9d .DUonjc .VfPpkd-LgbsSe:disabled.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:0;opacity:var(--mdc-ripple-hover-opacity,0)}.jR8x9d .DUonjc .VfPpkd-LgbsSe:disabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.jR8x9d .DUonjc .VfPpkd-LgbsSe:disabled:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:0;opacity:var(--mdc-ripple-focus-opacity,0)}.jR8x9d .DUonjc .VfPpkd-LgbsSe:disabled:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .DUonjc .VfPpkd-LgbsSe:disabled:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:0;opacity:var(--mdc-ripple-press-opacity,0)}.jR8x9d .DUonjc .VfPpkd-LgbsSe:disabled.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0)}.jR8x9d .DUonjc .UMrnmb-jsLfKf-JIbuQc{margin-right:8px}.jR8x9d .AjY5Oe{font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:.875rem;letter-spacing:.0107142857em;font-weight:500;text-transform:none;-webkit-transition:border .28s cubic-bezier(.4,0,.2,1),box-shadow .28s cubic-bezier(.4,0,.2,1);transition:border .28s cubic-bezier(.4,0,.2,1),box-shadow .28s cubic-bezier(.4,0,.2,1);box-shadow:none}.jR8x9d .AjY5Oe .VfPpkd-Jh9lGc{height:100%;position:absolute;overflow:hidden;width:100%;z-index:0}.jR8x9d .AjY5Oe:not(:disabled){background-color:rgb(138,180,248);background-color:var(--gm-fillbutton-container-color,rgb(138,180,248))}.jR8x9d .AjY5Oe:not(:disabled){color:rgb(32,33,36);color:var(--gm-fillbutton-ink-color,rgb(32,33,36))}.jR8x9d .AjY5Oe:disabled{background-color:rgba(232,234,237,.12);background-color:var(--gm-fillbutton-disabled-container-color,rgba(232,234,237,.12))}.jR8x9d .AjY5Oe:disabled{color:rgba(232,234,237,.38);color:var(--gm-fillbutton-disabled-ink-color,rgba(232,234,237,.38))}.jR8x9d .AjY5Oe .VfPpkd-Jh9lGc::before,.jR8x9d .AjY5Oe .VfPpkd-Jh9lGc::after{background-color:#fff;background-color:var(--gm-fillbutton-state-color,#fff)}.jR8x9d .AjY5Oe:hover .VfPpkd-Jh9lGc::before,.jR8x9d .AjY5Oe.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:.16;opacity:var(--mdc-ripple-hover-opacity,.16)}.jR8x9d .AjY5Oe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.jR8x9d .AjY5Oe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.24;opacity:var(--mdc-ripple-focus-opacity,.24)}.jR8x9d .AjY5Oe:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .AjY5Oe:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.2;opacity:var(--mdc-ripple-press-opacity,.2)}.jR8x9d .AjY5Oe.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.2)}.jR8x9d .AjY5Oe .VfPpkd-BFbNVe-bF1uUb{opacity:0}.jR8x9d .AjY5Oe .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo,.jR8x9d .AjY5Oe .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:rgb(32,33,36)}}@media screen and (prefers-color-scheme:dark) and (-ms-high-contrast:active),screen and (prefers-color-scheme:dark) and (forced-colors:active){.jR8x9d .AjY5Oe .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo,.jR8x9d .AjY5Oe .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:CanvasText}}@media screen and (prefers-color-scheme:dark){.jR8x9d .AjY5Oe:hover{box-shadow:0 1px 2px 0 rgba(0,0,0,.3),0 1px 3px 1px rgba(0,0,0,.15);box-shadow:0 1px 2px 0 var(--gm-fillbutton-keyshadow-color,rgba(0,0,0,.3)),0 1px 3px 1px var(--gm-fillbutton-ambientshadow-color,rgba(0,0,0,.15))}.jR8x9d .AjY5Oe:hover .VfPpkd-BFbNVe-bF1uUb{opacity:0}.jR8x9d .AjY5Oe:active{box-shadow:0 1px 2px 0 rgba(0,0,0,.3),0 2px 6px 2px rgba(0,0,0,.15);box-shadow:0 1px 2px 0 var(--gm-fillbutton-keyshadow-color,rgba(0,0,0,.3)),0 2px 6px 2px var(--gm-fillbutton-ambientshadow-color,rgba(0,0,0,.15))}.jR8x9d .AjY5Oe:active .VfPpkd-BFbNVe-bF1uUb{opacity:0}.jR8x9d .AjY5Oe:disabled{box-shadow:none}.jR8x9d .AjY5Oe:disabled:hover .VfPpkd-Jh9lGc::before,.jR8x9d .AjY5Oe:disabled.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:0;opacity:var(--mdc-ripple-hover-opacity,0)}.jR8x9d .AjY5Oe:disabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.jR8x9d .AjY5Oe:disabled:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:0;opacity:var(--mdc-ripple-focus-opacity,0)}.jR8x9d .AjY5Oe:disabled:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .AjY5Oe:disabled:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:0;opacity:var(--mdc-ripple-press-opacity,0)}.jR8x9d .AjY5Oe:disabled.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0)}.jR8x9d .AjY5Oe:disabled .VfPpkd-BFbNVe-bF1uUb{opacity:0}.jR8x9d .OLiIxf{font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:.875rem;letter-spacing:.0107142857em;font-weight:500;text-transform:none;-webkit-transition:border .28s cubic-bezier(.4,0,.2,1),box-shadow .28s cubic-bezier(.4,0,.2,1);transition:border .28s cubic-bezier(.4,0,.2,1),box-shadow .28s cubic-bezier(.4,0,.2,1);box-shadow:none}.jR8x9d .OLiIxf .VfPpkd-Jh9lGc{height:100%;position:absolute;overflow:hidden;width:100%;z-index:0}.jR8x9d .OLiIxf:not(:disabled){color:rgb(138,180,248);color:var(--gm-hairlinebutton-ink-color,rgb(138,180,248))}.jR8x9d .OLiIxf:not(:disabled){border-color:rgb(95,99,104);border-color:var(--gm-hairlinebutton-outline-color,rgb(95,99,104))}.jR8x9d .OLiIxf:not(:disabled):hover{border-color:rgb(95,99,104);border-color:var(--gm-hairlinebutton-outline-color,rgb(95,99,104))}.jR8x9d .OLiIxf:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.jR8x9d .OLiIxf:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{border-color:rgb(174,203,250);border-color:var(--gm-hairlinebutton-outline-color--stateful,rgb(174,203,250))}.jR8x9d .OLiIxf:not(:disabled):active,.jR8x9d .OLiIxf:not(:disabled):focus:active{border-color:rgb(95,99,104);border-color:var(--gm-hairlinebutton-outline-color,rgb(95,99,104))}.jR8x9d .OLiIxf:disabled{color:rgba(232,234,237,.38);color:var(--gm-hairlinebutton-disabled-ink-color,rgba(232,234,237,.38))}.jR8x9d .OLiIxf:disabled{border-color:rgba(232,234,237,.12);border-color:var(--gm-hairlinebutton-disabled-outline-color,rgba(232,234,237,.12))}.jR8x9d .OLiIxf:hover:not(:disabled),.jR8x9d .OLiIxf.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:disabled),.jR8x9d .OLiIxf:not(.VfPpkd-ksKsZd-mWPk3d):focus:not(:disabled),.jR8x9d .OLiIxf:active:not(:disabled){color:rgb(174,203,250);color:var(--gm-hairlinebutton-ink-color--stateful,rgb(174,203,250))}.jR8x9d .OLiIxf .VfPpkd-BFbNVe-bF1uUb{opacity:0}.jR8x9d .OLiIxf .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo,.jR8x9d .OLiIxf .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:rgb(138,180,248)}}@media screen and (prefers-color-scheme:dark) and (-ms-high-contrast:active),screen and (prefers-color-scheme:dark) and (forced-colors:active){.jR8x9d .OLiIxf .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo,.jR8x9d .OLiIxf .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:CanvasText}}@media screen and (prefers-color-scheme:dark){.jR8x9d .OLiIxf .VfPpkd-Jh9lGc::before,.jR8x9d .OLiIxf .VfPpkd-Jh9lGc::after{background-color:rgb(138,180,248);background-color:var(--gm-hairlinebutton-state-color,rgb(138,180,248))}.jR8x9d .OLiIxf:hover .VfPpkd-Jh9lGc::before,.jR8x9d .OLiIxf.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.jR8x9d .OLiIxf.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.jR8x9d .OLiIxf:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.jR8x9d .OLiIxf:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .OLiIxf:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.jR8x9d .OLiIxf.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}.jR8x9d .OLiIxf:disabled:hover .VfPpkd-Jh9lGc::before,.jR8x9d .OLiIxf:disabled.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:0;opacity:var(--mdc-ripple-hover-opacity,0)}.jR8x9d .OLiIxf:disabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.jR8x9d .OLiIxf:disabled:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:0;opacity:var(--mdc-ripple-focus-opacity,0)}.jR8x9d .OLiIxf:disabled:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .OLiIxf:disabled:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:0;opacity:var(--mdc-ripple-press-opacity,0)}.jR8x9d .OLiIxf:disabled.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0)}.jR8x9d .MQas1c{font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:.875rem;letter-spacing:.0107142857em;font-weight:500;text-transform:none;-webkit-transition:border .28s cubic-bezier(.4,0,.2,1),box-shadow .28s cubic-bezier(.4,0,.2,1);transition:border .28s cubic-bezier(.4,0,.2,1),box-shadow .28s cubic-bezier(.4,0,.2,1);border-width:0;box-shadow:0 1px 2px 0 rgba(0,0,0,.3),0 1px 3px 1px rgba(0,0,0,.15);box-shadow:0 1px 2px 0 var(--gm-protectedbutton-keyshadow-color,rgba(0,0,0,.3)),0 1px 3px 1px var(--gm-protectedbutton-ambientshadow-color,rgba(0,0,0,.15))}.jR8x9d .MQas1c .VfPpkd-Jh9lGc{height:100%;position:absolute;overflow:hidden;width:100%;z-index:0}.jR8x9d .MQas1c:not(:disabled){background-color:rgb(32,33,36);background-color:var(--gm-protectedbutton-container-color,rgb(32,33,36))}.jR8x9d .MQas1c:not(:disabled){color:rgb(138,180,248);color:var(--gm-protectedbutton-ink-color,rgb(138,180,248))}.jR8x9d .MQas1c:disabled{background-color:rgba(232,234,237,.12);background-color:var(--gm-protectedbutton-disabled-container-color,rgba(232,234,237,.12))}.jR8x9d .MQas1c:disabled{color:rgba(232,234,237,.38);color:var(--gm-protectedbutton-disabled-ink-color,rgba(232,234,237,.38))}.jR8x9d .MQas1c:hover:not(:disabled),.jR8x9d .MQas1c.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:disabled),.jR8x9d .MQas1c:not(.VfPpkd-ksKsZd-mWPk3d):focus:not(:disabled),.jR8x9d .MQas1c:active:not(:disabled){color:rgb(174,203,250);color:var(--gm-protectedbutton-ink-color--stateful,rgb(174,203,250))}.jR8x9d .MQas1c .VfPpkd-BFbNVe-bF1uUb{opacity:.05}.jR8x9d .MQas1c .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo,.jR8x9d .MQas1c .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:rgb(138,180,248)}}@media screen and (prefers-color-scheme:dark) and (-ms-high-contrast:active),screen and (prefers-color-scheme:dark) and (forced-colors:active){.jR8x9d .MQas1c .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo,.jR8x9d .MQas1c .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:CanvasText}}@media screen and (prefers-color-scheme:dark){.jR8x9d .MQas1c.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.jR8x9d .MQas1c:not(.VfPpkd-ksKsZd-mWPk3d):focus{border-width:0;box-shadow:0 1px 2px 0 rgba(0,0,0,.3),0 1px 3px 1px rgba(0,0,0,.15);box-shadow:0 1px 2px 0 var(--gm-protectedbutton-keyshadow-color,rgba(0,0,0,.3)),0 1px 3px 1px var(--gm-protectedbutton-ambientshadow-color,rgba(0,0,0,.15))}.jR8x9d .MQas1c.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-BFbNVe-bF1uUb,.jR8x9d .MQas1c:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-BFbNVe-bF1uUb{opacity:.05}.jR8x9d .MQas1c:hover{border-width:0;box-shadow:0 1px 2px 0 rgba(0,0,0,.3),0 2px 6px 2px rgba(0,0,0,.15);box-shadow:0 1px 2px 0 var(--gm-protectedbutton-keyshadow-color,rgba(0,0,0,.3)),0 2px 6px 2px var(--gm-protectedbutton-ambientshadow-color,rgba(0,0,0,.15))}.jR8x9d .MQas1c:hover .VfPpkd-BFbNVe-bF1uUb{opacity:.08}.jR8x9d .MQas1c:not(:disabled):active{border-width:0;box-shadow:0 1px 3px 0 rgba(0,0,0,.3),0 4px 8px 3px rgba(0,0,0,.15);box-shadow:0 1px 3px 0 var(--gm-protectedbutton-keyshadow-color,rgba(0,0,0,.3)),0 4px 8px 3px var(--gm-protectedbutton-ambientshadow-color,rgba(0,0,0,.15))}.jR8x9d .MQas1c:not(:disabled):active .VfPpkd-BFbNVe-bF1uUb{opacity:.11}.jR8x9d .MQas1c .VfPpkd-Jh9lGc::before,.jR8x9d .MQas1c .VfPpkd-Jh9lGc::after{background-color:rgb(174,203,250);background-color:var(--gm-protectedbutton-state-color,rgb(174,203,250))}.jR8x9d .MQas1c:hover .VfPpkd-Jh9lGc::before,.jR8x9d .MQas1c.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.jR8x9d .MQas1c.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.jR8x9d .MQas1c:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.jR8x9d .MQas1c:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .MQas1c:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.jR8x9d .MQas1c.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}.jR8x9d .MQas1c:disabled{border-width:0;box-shadow:0 1px 2px 0 rgba(0,0,0,.3),0 1px 3px 1px rgba(0,0,0,.15);box-shadow:0 1px 2px 0 var(--gm-protectedbutton-keyshadow-color,rgba(0,0,0,.3)),0 1px 3px 1px var(--gm-protectedbutton-ambientshadow-color,rgba(0,0,0,.15))}.jR8x9d .MQas1c:disabled .VfPpkd-BFbNVe-bF1uUb{opacity:.05}.jR8x9d .MQas1c:disabled:hover .VfPpkd-Jh9lGc::before,.jR8x9d .MQas1c:disabled.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:0;opacity:var(--mdc-ripple-hover-opacity,0)}.jR8x9d .MQas1c:disabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.jR8x9d .MQas1c:disabled:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:0;opacity:var(--mdc-ripple-focus-opacity,0)}.jR8x9d .MQas1c:disabled:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .MQas1c:disabled:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:0;opacity:var(--mdc-ripple-press-opacity,0)}.jR8x9d .MQas1c:disabled.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0)}.jR8x9d .C1Uh5b{font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:.875rem;letter-spacing:.0107142857em;font-weight:500;text-transform:none;-webkit-transition:border .28s cubic-bezier(.4,0,.2,1),box-shadow .28s cubic-bezier(.4,0,.2,1);transition:border .28s cubic-bezier(.4,0,.2,1),box-shadow .28s cubic-bezier(.4,0,.2,1);box-shadow:none}.jR8x9d .C1Uh5b .VfPpkd-Jh9lGc{height:100%;position:absolute;overflow:hidden;width:100%;z-index:0}.jR8x9d .C1Uh5b:not(:disabled){background-color:rgba(138,180,248,.24)}.jR8x9d .C1Uh5b:not(:disabled){color:rgb(210,227,252)}.jR8x9d .C1Uh5b:disabled{background-color:rgba(232,234,237,.12)}.jR8x9d .C1Uh5b:disabled{color:rgba(232,234,237,.38)}.jR8x9d .C1Uh5b:hover:not(:disabled),.jR8x9d .C1Uh5b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:disabled),.jR8x9d .C1Uh5b:not(.VfPpkd-ksKsZd-mWPk3d):focus:not(:disabled),.jR8x9d .C1Uh5b:active:not(:disabled){color:#fff}.jR8x9d .C1Uh5b .VfPpkd-Jh9lGc::before,.jR8x9d .C1Uh5b .VfPpkd-Jh9lGc::after{background-color:#fff;background-color:var(--mdc-ripple-color,#fff)}.jR8x9d .C1Uh5b:hover .VfPpkd-Jh9lGc::before,.jR8x9d .C1Uh5b.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.jR8x9d .C1Uh5b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.jR8x9d .C1Uh5b:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.jR8x9d .C1Uh5b:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .C1Uh5b:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.jR8x9d .C1Uh5b.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}.jR8x9d .C1Uh5b .VfPpkd-BFbNVe-bF1uUb{opacity:0}.jR8x9d .C1Uh5b .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo,.jR8x9d .C1Uh5b .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:rgb(210,227,252)}}@media screen and (prefers-color-scheme:dark) and (-ms-high-contrast:active),screen and (prefers-color-scheme:dark) and (forced-colors:active){.jR8x9d .C1Uh5b .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo,.jR8x9d .C1Uh5b .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:CanvasText}}@media screen and (prefers-color-scheme:dark){.jR8x9d .C1Uh5b:hover{box-shadow:0 1px 2px 0 rgba(0,0,0,.3),0 1px 3px 1px rgba(0,0,0,.15)}.jR8x9d .C1Uh5b:hover .VfPpkd-BFbNVe-bF1uUb{opacity:0}.jR8x9d .C1Uh5b:not(:disabled):active{box-shadow:0 1px 2px 0 rgba(0,0,0,.3),0 2px 6px 2px rgba(0,0,0,.15)}.jR8x9d .C1Uh5b:not(:disabled):active .VfPpkd-BFbNVe-bF1uUb{opacity:0}.jR8x9d .C1Uh5b:disabled{box-shadow:none}.jR8x9d .C1Uh5b:disabled .VfPpkd-BFbNVe-bF1uUb{opacity:0}.jR8x9d .C1Uh5b:disabled:hover .VfPpkd-Jh9lGc::before,.jR8x9d .C1Uh5b:disabled.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:0;opacity:var(--mdc-ripple-hover-opacity,0)}.jR8x9d .C1Uh5b:disabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.jR8x9d .C1Uh5b:disabled:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:0;opacity:var(--mdc-ripple-focus-opacity,0)}.jR8x9d .C1Uh5b:disabled:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .C1Uh5b:disabled:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:0;opacity:var(--mdc-ripple-press-opacity,0)}.jR8x9d .C1Uh5b:disabled.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0)}.jR8x9d .lKxP2d{font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:.875rem;letter-spacing:.0107142857em;font-weight:500;text-transform:none}.jR8x9d .lKxP2d .VfPpkd-Jh9lGc{height:100%;position:absolute;overflow:hidden;width:100%;z-index:0}.jR8x9d .lKxP2d:not(:disabled){background-color:transparent}.jR8x9d .lKxP2d:not(:disabled){color:rgb(138,180,248);color:var(--gm-colortextbutton-ink-color,rgb(138,180,248))}.jR8x9d .lKxP2d:disabled{color:rgba(232,234,237,.38);color:var(--gm-colortextbutton-disabled-ink-color,rgba(232,234,237,.38))}.jR8x9d .lKxP2d .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo,.jR8x9d .lKxP2d .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:rgb(138,180,248)}}@media screen and (prefers-color-scheme:dark) and (-ms-high-contrast:active),screen and (prefers-color-scheme:dark) and (forced-colors:active){.jR8x9d .lKxP2d .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo,.jR8x9d .lKxP2d .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:CanvasText}}@media screen and (prefers-color-scheme:dark){.jR8x9d .lKxP2d:hover:not(:disabled),.jR8x9d .lKxP2d.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:disabled),.jR8x9d .lKxP2d:not(.VfPpkd-ksKsZd-mWPk3d):focus:not(:disabled),.jR8x9d .lKxP2d:active:not(:disabled){color:rgb(174,203,250);color:var(--gm-colortextbutton-ink-color--stateful,rgb(174,203,250))}.jR8x9d .lKxP2d .VfPpkd-Jh9lGc::before,.jR8x9d .lKxP2d .VfPpkd-Jh9lGc::after{background-color:rgb(174,203,250);background-color:var(--gm-colortextbutton-state-color,rgb(174,203,250))}.jR8x9d .lKxP2d:hover .VfPpkd-Jh9lGc::before,.jR8x9d .lKxP2d.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.jR8x9d .lKxP2d.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.jR8x9d .lKxP2d:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.jR8x9d .lKxP2d:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .lKxP2d:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.jR8x9d .lKxP2d.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}.jR8x9d .lKxP2d:disabled:hover .VfPpkd-Jh9lGc::before,.jR8x9d .lKxP2d:disabled.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:0;opacity:var(--mdc-ripple-hover-opacity,0)}.jR8x9d .lKxP2d:disabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.jR8x9d .lKxP2d:disabled:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:0;opacity:var(--mdc-ripple-focus-opacity,0)}.jR8x9d .lKxP2d:disabled:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .lKxP2d:disabled:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:0;opacity:var(--mdc-ripple-press-opacity,0)}.jR8x9d .lKxP2d:disabled.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0)}.jR8x9d .XhPA0b{font-family:"Google Sans",Roboto,Arial,sans-serif;font-size:.875rem;letter-spacing:.0107142857em;font-weight:500;text-transform:none}.jR8x9d .XhPA0b .VfPpkd-Jh9lGc{height:100%;position:absolute;overflow:hidden;width:100%;z-index:0}.jR8x9d .XhPA0b:not(:disabled){color:rgb(232,234,237);color:var(--gm-neutraltextbutton-ink-color,rgb(232,234,237))}.jR8x9d .XhPA0b:disabled{color:rgba(232,234,237,.38);color:var(--gm-neutraltextbutton-disabled-ink-color,rgba(232,234,237,.38))}.jR8x9d .XhPA0b:hover:not(:disabled),.jR8x9d .XhPA0b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:disabled),.jR8x9d .XhPA0b:not(.VfPpkd-ksKsZd-mWPk3d):focus:not(:disabled),.jR8x9d .XhPA0b:active:not(:disabled){color:rgb(248,249,250);color:var(--gm-neutraltextbutton-ink-color--stateful,rgb(248,249,250))}.jR8x9d .XhPA0b .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo,.jR8x9d .XhPA0b .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:rgb(232,234,237)}}@media screen and (prefers-color-scheme:dark) and (-ms-high-contrast:active),screen and (prefers-color-scheme:dark) and (forced-colors:active){.jR8x9d .XhPA0b .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo,.jR8x9d .XhPA0b .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:CanvasText}}@media screen and (prefers-color-scheme:dark){.jR8x9d .XhPA0b .VfPpkd-Jh9lGc::before,.jR8x9d .XhPA0b .VfPpkd-Jh9lGc::after{background-color:rgb(232,234,237);background-color:var(--gm-neutraltextbutton-state-color,rgb(232,234,237))}.jR8x9d .XhPA0b:hover .VfPpkd-Jh9lGc::before,.jR8x9d .XhPA0b.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.jR8x9d .XhPA0b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.jR8x9d .XhPA0b:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.jR8x9d .XhPA0b:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .XhPA0b:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.jR8x9d .XhPA0b.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}.jR8x9d .XhPA0b:disabled:hover .VfPpkd-Jh9lGc::before,.jR8x9d .XhPA0b:disabled.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:0;opacity:var(--mdc-ripple-hover-opacity,0)}.jR8x9d .XhPA0b:disabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.jR8x9d .XhPA0b:disabled:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:0;opacity:var(--mdc-ripple-focus-opacity,0)}.jR8x9d .XhPA0b:disabled:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .XhPA0b:disabled:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:0;opacity:var(--mdc-ripple-press-opacity,0)}.jR8x9d .XhPA0b:disabled.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0)}.jR8x9d .eT1oJ{z-index:0}.jR8x9d .eT1oJ .VfPpkd-Bz112c-Jh9lGc::before,.jR8x9d .eT1oJ .VfPpkd-Bz112c-Jh9lGc::after{z-index:-1}.jR8x9d .eT1oJ:disabled{color:rgba(232,234,237,.38);color:var(--gm-iconbutton-disabled-ink-color,rgba(232,234,237,.38))}.jR8x9d .eT1oJ .VfPpkd-Bz112c-Jh9lGc::before,.jR8x9d .eT1oJ .VfPpkd-Bz112c-Jh9lGc::after{background-color:rgb(232,234,237);background-color:var(--mdc-ripple-color,rgb(232,234,237))}.jR8x9d .eT1oJ:hover .VfPpkd-Bz112c-Jh9lGc::before,.jR8x9d .eT1oJ.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Bz112c-Jh9lGc::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.jR8x9d .eT1oJ.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Bz112c-Jh9lGc::before,.jR8x9d .eT1oJ:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Bz112c-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.jR8x9d .eT1oJ:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Bz112c-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .eT1oJ:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Bz112c-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.jR8x9d .eT1oJ.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}.jR8x9d .eT1oJ:disabled:hover .VfPpkd-Jh9lGc::before,.jR8x9d .eT1oJ:disabled.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:0;opacity:var(--mdc-ripple-hover-opacity,0)}.jR8x9d .eT1oJ:disabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.jR8x9d .eT1oJ:disabled:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:0;opacity:var(--mdc-ripple-focus-opacity,0)}.jR8x9d .eT1oJ:disabled:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .eT1oJ:disabled:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:0;opacity:var(--mdc-ripple-press-opacity,0)}.jR8x9d .eT1oJ:disabled.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0)}.jR8x9d .tmJved{z-index:0}.jR8x9d .tmJved .VfPpkd-Bz112c-Jh9lGc::before,.jR8x9d .tmJved .VfPpkd-Bz112c-Jh9lGc::after{z-index:-1}.jR8x9d .tmJved:disabled{color:rgba(232,234,237,.38);color:var(--gm-iconbutton-disabled-ink-color,rgba(232,234,237,.38))}.jR8x9d .tmJved .VfPpkd-Bz112c-Jh9lGc::before,.jR8x9d .tmJved .VfPpkd-Bz112c-Jh9lGc::after{background-color:rgb(232,234,237);background-color:var(--mdc-ripple-color,rgb(232,234,237))}.jR8x9d .tmJved:hover .VfPpkd-Bz112c-Jh9lGc::before,.jR8x9d .tmJved.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Bz112c-Jh9lGc::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.jR8x9d .tmJved.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Bz112c-Jh9lGc::before,.jR8x9d .tmJved:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Bz112c-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.jR8x9d .tmJved:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Bz112c-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .tmJved:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Bz112c-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.jR8x9d .tmJved.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}.jR8x9d .tmJved:disabled:hover .VfPpkd-Jh9lGc::before,.jR8x9d .tmJved:disabled.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:0;opacity:var(--mdc-ripple-hover-opacity,0)}.jR8x9d .tmJved:disabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.jR8x9d .tmJved:disabled:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:0;opacity:var(--mdc-ripple-focus-opacity,0)}.jR8x9d .tmJved:disabled:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .tmJved:disabled:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:0;opacity:var(--mdc-ripple-press-opacity,0)}.jR8x9d .tmJved:disabled.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0)}.jR8x9d .AaN0Dd{background-color:rgb(32,33,36);border:1px solid rgb(95,99,104);box-shadow:none}.jR8x9d .AaN0Dd .VfPpkd-BFbNVe-bF1uUb{opacity:0}.jR8x9d .AaN0Dd .VfPpkd-EScbFb-JIbuQc .VfPpkd-FJ5hab::before,.jR8x9d .AaN0Dd .VfPpkd-EScbFb-JIbuQc .VfPpkd-FJ5hab::after{background-color:rgb(232,234,237);background-color:var(--mdc-ripple-color,rgb(232,234,237))}.jR8x9d .AaN0Dd .VfPpkd-EScbFb-JIbuQc:hover .VfPpkd-FJ5hab::before,.jR8x9d .AaN0Dd .VfPpkd-EScbFb-JIbuQc.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-FJ5hab::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.jR8x9d .AaN0Dd .VfPpkd-EScbFb-JIbuQc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-FJ5hab::before,.jR8x9d .AaN0Dd .VfPpkd-EScbFb-JIbuQc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-FJ5hab::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.jR8x9d .AaN0Dd .VfPpkd-EScbFb-JIbuQc:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-FJ5hab::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .AaN0Dd .VfPpkd-EScbFb-JIbuQc:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-FJ5hab::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.jR8x9d .AaN0Dd .VfPpkd-EScbFb-JIbuQc.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}.jR8x9d .AaN0Dd .VfPpkd-gBNGNe{z-index:1}.jR8x9d .BKdRne{background-color:rgb(32,33,36);border-width:0;box-shadow:0 1px 2px 0 rgba(0,0,0,.3),0 1px 3px 1px rgba(0,0,0,.15)}.jR8x9d .BKdRne .VfPpkd-BFbNVe-bF1uUb{opacity:.05}.jR8x9d .BKdRne .VfPpkd-EScbFb-JIbuQc .VfPpkd-FJ5hab::before,.jR8x9d .BKdRne .VfPpkd-EScbFb-JIbuQc .VfPpkd-FJ5hab::after{background-color:rgb(232,234,237);background-color:var(--mdc-ripple-color,rgb(232,234,237))}.jR8x9d .BKdRne .VfPpkd-EScbFb-JIbuQc:hover .VfPpkd-FJ5hab::before,.jR8x9d .BKdRne .VfPpkd-EScbFb-JIbuQc.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-FJ5hab::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.jR8x9d .BKdRne .VfPpkd-EScbFb-JIbuQc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-FJ5hab::before,.jR8x9d .BKdRne .VfPpkd-EScbFb-JIbuQc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-FJ5hab::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.jR8x9d .BKdRne .VfPpkd-EScbFb-JIbuQc:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-FJ5hab::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .BKdRne .VfPpkd-EScbFb-JIbuQc:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-FJ5hab::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.jR8x9d .BKdRne .VfPpkd-EScbFb-JIbuQc.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}.jR8x9d .BKdRne .VfPpkd-gBNGNe{z-index:1}.jR8x9d .swXlm .VfPpkd-muHVFf-bMcfAe[disabled]:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:rgba(232,234,237,.38);border-color:var(--mdc-checkbox-disabled-unselected-icon-color,rgba(232,234,237,.38));background-color:transparent}.jR8x9d .swXlm .VfPpkd-muHVFf-bMcfAe[disabled]:checked~.VfPpkd-YQoJzd,.jR8x9d .swXlm .VfPpkd-muHVFf-bMcfAe[disabled]:indeterminate~.VfPpkd-YQoJzd,.jR8x9d .swXlm .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true][disabled]~.VfPpkd-YQoJzd{border-color:transparent;background-color:rgba(232,234,237,.38);background-color:var(--mdc-checkbox-disabled-selected-icon-color,rgba(232,234,237,.38))}.jR8x9d .swXlm .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd .VfPpkd-HUofsb{color:#202124;color:var(--mdc-checkbox-selected-checkmark-color,#202124)}.jR8x9d .swXlm .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd .VfPpkd-SJnn3d{border-color:#202124;border-color:var(--mdc-checkbox-selected-checkmark-color,#202124)}.jR8x9d .swXlm .VfPpkd-muHVFf-bMcfAe:disabled~.VfPpkd-YQoJzd .VfPpkd-HUofsb{color:#202124;color:var(--mdc-checkbox-disabled-selected-checkmark-color,#202124)}.jR8x9d .swXlm .VfPpkd-muHVFf-bMcfAe:disabled~.VfPpkd-YQoJzd .VfPpkd-SJnn3d{border-color:#202124;border-color:var(--mdc-checkbox-disabled-selected-checkmark-color,#202124)}.jR8x9d .swXlm .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:#9aa0a6;border-color:var(--mdc-checkbox-unselected-icon-color,#9aa0a6);background-color:transparent}.jR8x9d .swXlm .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.jR8x9d .swXlm .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.jR8x9d .swXlm .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd{border-color:#8ab4f8;border-color:var(--mdc-checkbox-selected-icon-color,#8ab4f8);background-color:#8ab4f8;background-color:var(--mdc-checkbox-selected-icon-color,#8ab4f8)}@-webkit-keyframes mdc-checkbox-fade-in-background-FF9AA0A6FF8AB4F800000000FF8AB4F8{0%{border-color:#9aa0a6;border-color:var(--mdc-checkbox-unselected-icon-color,#9aa0a6);background-color:transparent}50%{border-color:#8ab4f8;border-color:var(--mdc-checkbox-selected-icon-color,#8ab4f8);background-color:#8ab4f8;background-color:var(--mdc-checkbox-selected-icon-color,#8ab4f8)}}@keyframes mdc-checkbox-fade-in-background-FF9AA0A6FF8AB4F800000000FF8AB4F8{0%{border-color:#9aa0a6;border-color:var(--mdc-checkbox-unselected-icon-color,#9aa0a6);background-color:transparent}50%{border-color:#8ab4f8;border-color:var(--mdc-checkbox-selected-icon-color,#8ab4f8);background-color:#8ab4f8;background-color:var(--mdc-checkbox-selected-icon-color,#8ab4f8)}}@-webkit-keyframes mdc-checkbox-fade-out-background-FF9AA0A6FF8AB4F800000000FF8AB4F8{0%,80%{border-color:#8ab4f8;border-color:var(--mdc-checkbox-selected-icon-color,#8ab4f8);background-color:#8ab4f8;background-color:var(--mdc-checkbox-selected-icon-color,#8ab4f8)}100%{border-color:#9aa0a6;border-color:var(--mdc-checkbox-unselected-icon-color,#9aa0a6);background-color:transparent}}@keyframes mdc-checkbox-fade-out-background-FF9AA0A6FF8AB4F800000000FF8AB4F8{0%,80%{border-color:#8ab4f8;border-color:var(--mdc-checkbox-selected-icon-color,#8ab4f8);background-color:#8ab4f8;background-color:var(--mdc-checkbox-selected-icon-color,#8ab4f8)}100%{border-color:#9aa0a6;border-color:var(--mdc-checkbox-unselected-icon-color,#9aa0a6);background-color:transparent}}.jR8x9d .swXlm.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.jR8x9d .swXlm.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{-webkit-animation-name:mdc-checkbox-fade-in-background-FF9AA0A6FF8AB4F800000000FF8AB4F8;animation-name:mdc-checkbox-fade-in-background-FF9AA0A6FF8AB4F800000000FF8AB4F8}.jR8x9d .swXlm.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.jR8x9d .swXlm.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{-webkit-animation-name:mdc-checkbox-fade-out-background-FF9AA0A6FF8AB4F800000000FF8AB4F8;animation-name:mdc-checkbox-fade-out-background-FF9AA0A6FF8AB4F800000000FF8AB4F8}.jR8x9d .swXlm:hover .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:#f8f9fa;border-color:var(--mdc-checkbox-unselected-hover-icon-color,#f8f9fa);background-color:transparent}.jR8x9d .swXlm:hover .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.jR8x9d .swXlm:hover .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.jR8x9d .swXlm:hover .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd{border-color:#aecbfa;border-color:var(--mdc-checkbox-selected-hover-icon-color,#aecbfa);background-color:#aecbfa;background-color:var(--mdc-checkbox-selected-hover-icon-color,#aecbfa)}@-webkit-keyframes mdc-checkbox-fade-in-background-FFF8F9FAFFAECBFA00000000FFAECBFA{0%{border-color:#f8f9fa;border-color:var(--mdc-checkbox-unselected-hover-icon-color,#f8f9fa);background-color:transparent}50%{border-color:#aecbfa;border-color:var(--mdc-checkbox-selected-hover-icon-color,#aecbfa);background-color:#aecbfa;background-color:var(--mdc-checkbox-selected-hover-icon-color,#aecbfa)}}@-webkit-keyframes mdc-checkbox-fade-out-background-FFF8F9FAFFAECBFA00000000FFAECBFA{0%,80%{border-color:#aecbfa;border-color:var(--mdc-checkbox-selected-hover-icon-color,#aecbfa);background-color:#aecbfa;background-color:var(--mdc-checkbox-selected-hover-icon-color,#aecbfa)}100%{border-color:#f8f9fa;border-color:var(--mdc-checkbox-unselected-hover-icon-color,#f8f9fa);background-color:transparent}}.jR8x9d .swXlm:hover.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.jR8x9d .swXlm:hover.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{-webkit-animation-name:mdc-checkbox-fade-in-background-FFF8F9FAFFAECBFA00000000FFAECBFA;animation-name:mdc-checkbox-fade-in-background-FFF8F9FAFFAECBFA00000000FFAECBFA}.jR8x9d .swXlm:hover.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.jR8x9d .swXlm:hover.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{-webkit-animation-name:mdc-checkbox-fade-out-background-FFF8F9FAFFAECBFA00000000FFAECBFA;animation-name:mdc-checkbox-fade-out-background-FFF8F9FAFFAECBFA00000000FFAECBFA}.jR8x9d .swXlm.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd,.jR8x9d .swXlm:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:#f8f9fa;border-color:var(--mdc-checkbox-unselected-focus-icon-color,#f8f9fa);background-color:transparent}.jR8x9d .swXlm.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.jR8x9d .swXlm.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.jR8x9d .swXlm.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd,.jR8x9d .swXlm:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.jR8x9d .swXlm:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.jR8x9d .swXlm:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd{border-color:#aecbfa;border-color:var(--mdc-checkbox-selected-focus-icon-color,#aecbfa);background-color:#aecbfa;background-color:var(--mdc-checkbox-selected-focus-icon-color,#aecbfa)}.jR8x9d .swXlm.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.jR8x9d .swXlm.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.jR8x9d .swXlm:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.jR8x9d .swXlm:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{-webkit-animation-name:mdc-checkbox-fade-in-background-FFF8F9FAFFAECBFA00000000FFAECBFA;animation-name:mdc-checkbox-fade-in-background-FFF8F9FAFFAECBFA00000000FFAECBFA}.jR8x9d .swXlm.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.jR8x9d .swXlm.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.jR8x9d .swXlm:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.jR8x9d .swXlm:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{-webkit-animation-name:mdc-checkbox-fade-out-background-FFF8F9FAFFAECBFA00000000FFAECBFA;animation-name:mdc-checkbox-fade-out-background-FFF8F9FAFFAECBFA00000000FFAECBFA}.jR8x9d .swXlm:not(:disabled):active .VfPpkd-muHVFf-bMcfAe:enabled:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:#f8f9fa;border-color:var(--mdc-checkbox-unselected-pressed-icon-color,#f8f9fa);background-color:transparent}.jR8x9d .swXlm:not(:disabled):active .VfPpkd-muHVFf-bMcfAe:enabled:checked~.VfPpkd-YQoJzd,.jR8x9d .swXlm:not(:disabled):active .VfPpkd-muHVFf-bMcfAe:enabled:indeterminate~.VfPpkd-YQoJzd,.jR8x9d .swXlm:not(:disabled):active .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true]:enabled~.VfPpkd-YQoJzd{border-color:#aecbfa;border-color:var(--mdc-checkbox-selected-pressed-icon-color,#aecbfa);background-color:#aecbfa;background-color:var(--mdc-checkbox-selected-pressed-icon-color,#aecbfa)}@keyframes mdc-checkbox-fade-in-background-FFF8F9FAFFAECBFA00000000FFAECBFA{0%{border-color:#f8f9fa;border-color:var(--mdc-checkbox-unselected-pressed-icon-color,#f8f9fa);background-color:transparent}50%{border-color:#aecbfa;border-color:var(--mdc-checkbox-selected-pressed-icon-color,#aecbfa);background-color:#aecbfa;background-color:var(--mdc-checkbox-selected-pressed-icon-color,#aecbfa)}}@keyframes mdc-checkbox-fade-out-background-FFF8F9FAFFAECBFA00000000FFAECBFA{0%,80%{border-color:#aecbfa;border-color:var(--mdc-checkbox-selected-pressed-icon-color,#aecbfa);background-color:#aecbfa;background-color:var(--mdc-checkbox-selected-pressed-icon-color,#aecbfa)}100%{border-color:#f8f9fa;border-color:var(--mdc-checkbox-unselected-pressed-icon-color,#f8f9fa);background-color:transparent}}.jR8x9d .swXlm:not(:disabled):active.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-barxie .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.jR8x9d .swXlm:not(:disabled):active.VfPpkd-MPu53c-OWXEXe-vwu2ne-iAfbIe-A9y3zc .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{-webkit-animation-name:mdc-checkbox-fade-in-background-FFF8F9FAFFAECBFA00000000FFAECBFA;animation-name:mdc-checkbox-fade-in-background-FFF8F9FAFFAECBFA00000000FFAECBFA}.jR8x9d .swXlm:not(:disabled):active.VfPpkd-MPu53c-OWXEXe-vwu2ne-barxie-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd,.jR8x9d .swXlm:not(:disabled):active.VfPpkd-MPu53c-OWXEXe-vwu2ne-A9y3zc-iAfbIe .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd{-webkit-animation-name:mdc-checkbox-fade-out-background-FFF8F9FAFFAECBFA00000000FFAECBFA;animation-name:mdc-checkbox-fade-out-background-FFF8F9FAFFAECBFA00000000FFAECBFA}.jR8x9d .swXlm .VfPpkd-OYHm6b::before,.jR8x9d .swXlm .VfPpkd-OYHm6b::after{background-color:#e8eaed;background-color:var(--mdc-checkbox-unselected-hover-state-layer-color,#e8eaed)}.jR8x9d .swXlm:hover .VfPpkd-OYHm6b::before,.jR8x9d .swXlm.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-OYHm6b::before{opacity:.04;opacity:var(--mdc-checkbox-unselected-hover-state-layer-opacity,.04)}.jR8x9d .swXlm.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-OYHm6b::before,.jR8x9d .swXlm:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-OYHm6b::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-checkbox-unselected-focus-state-layer-opacity,.12)}.jR8x9d .swXlm:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-OYHm6b::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .swXlm:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-OYHm6b::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-checkbox-unselected-pressed-state-layer-opacity,.1)}.jR8x9d .swXlm.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-checkbox-unselected-pressed-state-layer-opacity,0.1)}.jR8x9d .swXlm .VfPpkd-OYHm6b::before{background-color:#e8eaed;background-color:var(--mdc-checkbox-unselected-hover-state-layer-color,#e8eaed)}.jR8x9d .swXlm .VfPpkd-OYHm6b::after{background-color:#8ab4f8;background-color:var(--mdc-checkbox-unselected-pressed-state-layer-color,#8ab4f8)}.jR8x9d .swXlm.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::before,.jR8x9d .swXlm.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::after{background-color:#8ab4f8;background-color:var(--mdc-checkbox-selected-hover-state-layer-color,#8ab4f8)}.jR8x9d .swXlm.VfPpkd-MPu53c-OWXEXe-gk6SMd:hover .VfPpkd-OYHm6b::before,.jR8x9d .swXlm.VfPpkd-MPu53c-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-OYHm6b::before{opacity:.04;opacity:var(--mdc-checkbox-selected-hover-state-layer-opacity,.04)}.jR8x9d .swXlm.VfPpkd-MPu53c-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-OYHm6b::before,.jR8x9d .swXlm.VfPpkd-MPu53c-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-OYHm6b::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-checkbox-selected-focus-state-layer-opacity,.12)}.jR8x9d .swXlm.VfPpkd-MPu53c-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-OYHm6b::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .swXlm.VfPpkd-MPu53c-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-OYHm6b::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-checkbox-selected-pressed-state-layer-opacity,.1)}.jR8x9d .swXlm.VfPpkd-MPu53c-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-checkbox-selected-pressed-state-layer-opacity,0.1)}.jR8x9d .swXlm.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::before,.jR8x9d .swXlm.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-MPu53c-OWXEXe-gk6SMd .VfPpkd-OYHm6b::after{background-color:#8ab4f8;background-color:var(--mdc-checkbox-selected-hover-state-layer-color,#8ab4f8)}}@media screen and (prefers-color-scheme:dark) and (forced-colors:active){.jR8x9d .swXlm .VfPpkd-muHVFf-bMcfAe[disabled]:not(:checked):not(:indeterminate):not([data-indeterminate=true])~.VfPpkd-YQoJzd{border-color:GrayText;border-color:var(--mdc-checkbox-disabled-unselected-icon-color,GrayText);background-color:transparent}.jR8x9d .swXlm .VfPpkd-muHVFf-bMcfAe[disabled]:checked~.VfPpkd-YQoJzd,.jR8x9d .swXlm .VfPpkd-muHVFf-bMcfAe[disabled]:indeterminate~.VfPpkd-YQoJzd,.jR8x9d .swXlm .VfPpkd-muHVFf-bMcfAe[data-indeterminate=true][disabled]~.VfPpkd-YQoJzd{border-color:GrayText;background-color:GrayText;background-color:var(--mdc-checkbox-disabled-selected-icon-color,GrayText)}.jR8x9d .swXlm .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd .VfPpkd-HUofsb{color:ButtonText;color:var(--mdc-checkbox-selected-checkmark-color,ButtonText)}.jR8x9d .swXlm .VfPpkd-muHVFf-bMcfAe:enabled~.VfPpkd-YQoJzd .VfPpkd-SJnn3d{border-color:ButtonText;border-color:var(--mdc-checkbox-selected-checkmark-color,ButtonText)}.jR8x9d .swXlm .VfPpkd-muHVFf-bMcfAe:disabled~.VfPpkd-YQoJzd .VfPpkd-HUofsb{color:ButtonFace;color:var(--mdc-checkbox-disabled-selected-checkmark-color,ButtonFace)}.jR8x9d .swXlm .VfPpkd-muHVFf-bMcfAe:disabled~.VfPpkd-YQoJzd .VfPpkd-SJnn3d{border-color:ButtonFace;border-color:var(--mdc-checkbox-disabled-selected-checkmark-color,ButtonFace)}}@media screen and (prefers-color-scheme:dark){.jR8x9d .MhRzze{font-family:"Google Sans",Roboto,Arial,sans-serif;line-height:1.25rem;font-size:.875rem;letter-spacing:.0178571429em;font-weight:500;-webkit-transition:box-shadow .28s cubic-bezier(.4,0,.2,1);transition:box-shadow .28s cubic-bezier(.4,0,.2,1);z-index:0;color:rgb(154,160,166);color:var(--gm-chip-ink-color,rgb(154,160,166))}.jR8x9d .MhRzze.VfPpkd-XPtOyb-OWXEXe-SNIJTd{-webkit-transition:box-shadow .28s cubic-bezier(.4,0,.2,1),opacity 75ms cubic-bezier(.4,0,.2,1),width .15s cubic-bezier(0,0,.2,1),padding .1s linear,margin .1s linear;transition:box-shadow .28s cubic-bezier(.4,0,.2,1),opacity 75ms cubic-bezier(.4,0,.2,1),width .15s cubic-bezier(0,0,.2,1),padding .1s linear,margin .1s linear}.jR8x9d .MhRzze .VfPpkd-v1cqY::before,.jR8x9d .MhRzze .VfPpkd-v1cqY::after{z-index:-1}.jR8x9d .MhRzze .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc{color:#9aa0a6}.jR8x9d .MhRzze .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc{color:rgb(154,160,166);color:var(--gm-chip-ink-color,rgb(154,160,166))}.jR8x9d .MhRzze .VfPpkd-Zr1Nwf-OWXEXe-UbuQg{color:#9aa0a6}.jR8x9d .MhRzze .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:hover{color:#9aa0a6}.jR8x9d .MhRzze .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:focus{color:#9aa0a6}.jR8x9d .MhRzze .VfPpkd-PvL5qd-Jt5cK{stroke:rgb(154,160,166);stroke:var(--gm-chip-ink-color,rgb(154,160,166))}.jR8x9d .MhRzze:hover,.jR8x9d .MhRzze.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.jR8x9d .MhRzze:not(.VfPpkd-ksKsZd-mWPk3d):focus,.jR8x9d .MhRzze:active{color:rgb(232,234,237);color:var(--gm-chip-ink-color--stateful,rgb(232,234,237))}.jR8x9d .MhRzze:hover .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc,.jR8x9d .MhRzze.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc,.jR8x9d .MhRzze:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc,.jR8x9d .MhRzze:active .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc{color:#e8eaed}.jR8x9d .MhRzze:hover .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc,.jR8x9d .MhRzze.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc,.jR8x9d .MhRzze:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc,.jR8x9d .MhRzze:active .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc{color:rgb(232,234,237);color:var(--gm-chip-ink-color--stateful,rgb(232,234,237))}.jR8x9d .MhRzze:hover .VfPpkd-Zr1Nwf-OWXEXe-UbuQg,.jR8x9d .MhRzze.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Zr1Nwf-OWXEXe-UbuQg,.jR8x9d .MhRzze:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Zr1Nwf-OWXEXe-UbuQg,.jR8x9d .MhRzze:active .VfPpkd-Zr1Nwf-OWXEXe-UbuQg{color:#e8eaed}.jR8x9d .MhRzze:hover .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:hover,.jR8x9d .MhRzze.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:hover,.jR8x9d .MhRzze:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:hover,.jR8x9d .MhRzze:active .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:hover{color:#e8eaed}.jR8x9d .MhRzze:hover .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:focus,.jR8x9d .MhRzze.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:focus,.jR8x9d .MhRzze:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:focus,.jR8x9d .MhRzze:active .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:focus{color:#e8eaed}.jR8x9d .MhRzze:hover .VfPpkd-PvL5qd-Jt5cK,.jR8x9d .MhRzze.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-PvL5qd-Jt5cK,.jR8x9d .MhRzze:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-PvL5qd-Jt5cK,.jR8x9d .MhRzze:active .VfPpkd-PvL5qd-Jt5cK{stroke:rgb(232,234,237);stroke:var(--gm-chip-ink-color--stateful,rgb(232,234,237))}.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd{background-color:rgba(138,180,248,.24);background-color:var(--gm-chip-container-color,rgba(138,180,248,.24));color:rgb(210,227,252);color:var(--gm-chip-ink-color,rgb(210,227,252));border-color:transparent;border-color:var(--gm-chip-outline-color--stateful,transparent)}.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc{color:#d2e3fc}.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc{color:rgb(210,227,252);color:var(--gm-chip-ink-color,rgb(210,227,252))}.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-Zr1Nwf-OWXEXe-UbuQg{color:#d2e3fc}.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:hover{color:#d2e3fc}.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:focus{color:#d2e3fc}.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-PvL5qd-Jt5cK{stroke:rgb(210,227,252);stroke:var(--gm-chip-ink-color,rgb(210,227,252))}.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd:hover,.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus,.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd:active{color:#fff;color:var(--gm-chip-ink-color--stateful,#fff)}.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd:hover .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc,.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc,.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc,.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd:active .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc{color:white}.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd:hover .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc,.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc,.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc,.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd:active .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc{color:#fff;color:var(--gm-chip-ink-color--stateful,#fff)}.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd:hover .VfPpkd-Zr1Nwf-OWXEXe-UbuQg,.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Zr1Nwf-OWXEXe-UbuQg,.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Zr1Nwf-OWXEXe-UbuQg,.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd:active .VfPpkd-Zr1Nwf-OWXEXe-UbuQg{color:white}.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd:hover .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:hover,.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:hover,.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:hover,.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd:active .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:hover{color:white}.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd:hover .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:focus,.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:focus,.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:focus,.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd:active .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:focus{color:white}.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd:hover .VfPpkd-PvL5qd-Jt5cK,.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-PvL5qd-Jt5cK,.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-PvL5qd-Jt5cK,.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd:active .VfPpkd-PvL5qd-Jt5cK{stroke:#fff;stroke:var(--gm-chip-ink-color--stateful,#fff)}.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-BFbNVe-bF1uUb{opacity:0}.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-v1cqY::before,.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-v1cqY::after{background-color:rgb(210,227,252);background-color:var(--gm-chip-state-color,rgb(210,227,252))}.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd:hover .VfPpkd-v1cqY::before,.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-v1cqY::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-v1cqY::before,.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-v1cqY::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-v1cqY::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-v1cqY::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.jR8x9d .MhRzze.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}.jR8x9d .fNK4Mb{background-color:rgb(32,33,36);background-color:var(--gm-chip-container-color,rgb(32,33,36));padding-right:16px;padding-left:16px;border-width:0;box-shadow:0 1px 2px 0 rgba(0,0,0,.3),0 1px 3px 1px rgba(0,0,0,.15)}.jR8x9d .fNK4Mb .VfPpkd-v1cqY::before,.jR8x9d .fNK4Mb .VfPpkd-v1cqY::after{background-color:rgb(232,234,237);background-color:var(--gm-chip-state-color,rgb(232,234,237))}.jR8x9d .fNK4Mb:hover .VfPpkd-v1cqY::before,.jR8x9d .fNK4Mb.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-v1cqY::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.jR8x9d .fNK4Mb.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-v1cqY::before,.jR8x9d .fNK4Mb:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-v1cqY::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.jR8x9d .fNK4Mb:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-v1cqY::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .fNK4Mb:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-v1cqY::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.jR8x9d .fNK4Mb.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}.jR8x9d .fNK4Mb .VfPpkd-BFbNVe-bF1uUb{opacity:.05}.jR8x9d .fNK4Mb:hover{border-width:0;box-shadow:0 1px 2px 0 rgba(0,0,0,.3),0 2px 6px 2px rgba(0,0,0,.15)}.jR8x9d .fNK4Mb:hover .VfPpkd-BFbNVe-bF1uUb{opacity:.08}.jR8x9d .fNK4Mb:active{border-width:0;box-shadow:0 1px 3px 0 rgba(0,0,0,.3),0 4px 8px 3px rgba(0,0,0,.15)}.jR8x9d .fNK4Mb:active .VfPpkd-BFbNVe-bF1uUb{opacity:.11}.jR8x9d .EuHQ0d{background-color:transparent;background-color:var(--gm-chip-container-color,transparent);border-style:solid;padding-right:15px;padding-left:15px;border-width:1px;border-color:rgb(95,99,104);border-color:var(--gm-chip-outline-color,rgb(95,99,104))}.jR8x9d .EuHQ0d .VfPpkd-v1cqY{top:-1px;left:-1px;border:1px solid transparent}.jR8x9d .EuHQ0d .VfPpkd-v1cqY::before,.jR8x9d .EuHQ0d .VfPpkd-v1cqY::after{background-color:rgb(232,234,237);background-color:var(--gm-chip-state-color,rgb(232,234,237))}.jR8x9d .EuHQ0d:hover .VfPpkd-v1cqY::before,.jR8x9d .EuHQ0d.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-v1cqY::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.jR8x9d .EuHQ0d.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-v1cqY::before,.jR8x9d .EuHQ0d:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-v1cqY::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.jR8x9d .EuHQ0d:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-v1cqY::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .EuHQ0d:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-v1cqY::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.jR8x9d .EuHQ0d.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}.jR8x9d .EuHQ0d:focus,.jR8x9d .EuHQ0d.VfPpkd-XPtOyb-OWXEXe-ssJRIf-JIbuQc-XpnDCe{border-color:rgb(232,234,237);border-color:var(--gm-chip-outline-color--stateful,rgb(232,234,237))}.jR8x9d .EuHQ0d:active{box-shadow:none}.jR8x9d .EuHQ0d:active .VfPpkd-BFbNVe-bF1uUb{opacity:0}.jR8x9d .EuHQ0d.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd{padding-right:16px;padding-left:16px;border-width:0}.jR8x9d .EuHQ0d.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-v1cqY{top:0;left:0;border:0 solid transparent}.jR8x9d .EuHQ0d.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd:hover{box-shadow:0 1px 2px 0 rgba(0,0,0,.3),0 1px 3px 1px rgba(0,0,0,.15)}.jR8x9d .EuHQ0d.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd:hover .VfPpkd-BFbNVe-bF1uUb{opacity:0}.jR8x9d .EuHQ0d.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd:focus,.jR8x9d .EuHQ0d.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd.VfPpkd-XPtOyb-OWXEXe-ssJRIf-JIbuQc-XpnDCe{padding-right:15px;padding-left:15px;border-width:1px}.jR8x9d .EuHQ0d.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd:focus .VfPpkd-v1cqY,.jR8x9d .EuHQ0d.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd.VfPpkd-XPtOyb-OWXEXe-ssJRIf-JIbuQc-XpnDCe .VfPpkd-v1cqY{top:-1px;left:-1px;border:1px solid transparent}.jR8x9d .X4PEqe{color:rgb(232,234,237);color:var(--gm-chip-ink-color,rgb(232,234,237))}.jR8x9d .X4PEqe .VfPpkd-Zr1Nwf.VfPpkd-Zr1Nwf-OWXEXe-M1Soyc:not(.VfPpkd-Zr1Nwf-OWXEXe-M1Soyc-L6cTce){width:20px;height:20px;font-size:20px}.jR8x9d .X4PEqe.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-PvL5qd,.jR8x9d .X4PEqe .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc:not(.VfPpkd-Zr1Nwf-OWXEXe-M1Soyc-L6cTce){margin-left:-8px;margin-right:8px}[dir=rtl] .jR8x9d .X4PEqe.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-PvL5qd,[dir=rtl] .jR8x9d .X4PEqe .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc:not(.VfPpkd-Zr1Nwf-OWXEXe-M1Soyc-L6cTce),.jR8x9d .X4PEqe.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-PvL5qd[dir=rtl],.jR8x9d .X4PEqe .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc:not(.VfPpkd-Zr1Nwf-OWXEXe-M1Soyc-L6cTce)[dir=rtl]{margin-left:8px;margin-right:-8px}.jR8x9d .X4PEqe .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc{color:#e8eaed}.jR8x9d .X4PEqe .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc{color:rgb(232,234,237);color:var(--gm-chip-ink-color,rgb(232,234,237))}.jR8x9d .X4PEqe .VfPpkd-Zr1Nwf-OWXEXe-UbuQg{color:#e8eaed}.jR8x9d .X4PEqe .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:hover{color:#e8eaed}.jR8x9d .X4PEqe .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:focus{color:#e8eaed}.jR8x9d .X4PEqe .VfPpkd-PvL5qd-Jt5cK{stroke:rgb(232,234,237);stroke:var(--gm-chip-ink-color,rgb(232,234,237))}.jR8x9d .X4PEqe:hover,.jR8x9d .X4PEqe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.jR8x9d .X4PEqe:not(.VfPpkd-ksKsZd-mWPk3d):focus,.jR8x9d .X4PEqe:active{color:rgb(248,249,250);color:var(--gm-chip-ink-color--stateful,rgb(248,249,250))}.jR8x9d .X4PEqe:hover .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc,.jR8x9d .X4PEqe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc,.jR8x9d .X4PEqe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc,.jR8x9d .X4PEqe:active .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc{color:#f8f9fa}.jR8x9d .X4PEqe:hover .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc,.jR8x9d .X4PEqe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc,.jR8x9d .X4PEqe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc,.jR8x9d .X4PEqe:active .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc{color:rgb(248,249,250);color:var(--gm-chip-ink-color--stateful,rgb(248,249,250))}.jR8x9d .X4PEqe:hover .VfPpkd-Zr1Nwf-OWXEXe-UbuQg,.jR8x9d .X4PEqe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Zr1Nwf-OWXEXe-UbuQg,.jR8x9d .X4PEqe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Zr1Nwf-OWXEXe-UbuQg,.jR8x9d .X4PEqe:active .VfPpkd-Zr1Nwf-OWXEXe-UbuQg{color:#f8f9fa}.jR8x9d .X4PEqe:hover .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:hover,.jR8x9d .X4PEqe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:hover,.jR8x9d .X4PEqe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:hover,.jR8x9d .X4PEqe:active .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:hover{color:#f8f9fa}.jR8x9d .X4PEqe:hover .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:focus,.jR8x9d .X4PEqe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:focus,.jR8x9d .X4PEqe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:focus,.jR8x9d .X4PEqe:active .VfPpkd-Zr1Nwf-OWXEXe-UbuQg:focus{color:#f8f9fa}.jR8x9d .X4PEqe:hover .VfPpkd-PvL5qd-Jt5cK,.jR8x9d .X4PEqe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-PvL5qd-Jt5cK,.jR8x9d .X4PEqe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-PvL5qd-Jt5cK,.jR8x9d .X4PEqe:active .VfPpkd-PvL5qd-Jt5cK{stroke:rgb(248,249,250);stroke:var(--gm-chip-ink-color--stateful,rgb(248,249,250))}.jR8x9d .Vo0FCd{font-family:Roboto,Arial,sans-serif;line-height:1.25rem;font-size:.875rem;letter-spacing:.0178571429em;font-weight:500;padding-right:11px;padding-left:11px;border-width:1px}.jR8x9d .Vo0FCd .VfPpkd-Zr1Nwf.VfPpkd-Zr1Nwf-OWXEXe-M1Soyc:not(.VfPpkd-Zr1Nwf-OWXEXe-M1Soyc-L6cTce){width:20px;height:20px;font-size:20px}.jR8x9d .Vo0FCd.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-PvL5qd,.jR8x9d .Vo0FCd .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc:not(.VfPpkd-Zr1Nwf-OWXEXe-M1Soyc-L6cTce){margin-left:-3px;margin-right:8px}[dir=rtl] .jR8x9d .Vo0FCd.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-PvL5qd,[dir=rtl] .jR8x9d .Vo0FCd .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc:not(.VfPpkd-Zr1Nwf-OWXEXe-M1Soyc-L6cTce),.jR8x9d .Vo0FCd.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-PvL5qd[dir=rtl],.jR8x9d .Vo0FCd .VfPpkd-Zr1Nwf-OWXEXe-M1Soyc:not(.VfPpkd-Zr1Nwf-OWXEXe-M1Soyc-L6cTce)[dir=rtl]{margin-left:8px;margin-right:-3px}.jR8x9d .Vo0FCd .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc{margin-left:8px;margin-right:-7px}[dir=rtl] .jR8x9d .Vo0FCd .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc,.jR8x9d .Vo0FCd .VfPpkd-StrnGf-XPtOyb-UbuQg-JIbuQc[dir=rtl]{margin-left:-7px;margin-right:8px}.jR8x9d .Vo0FCd .VfPpkd-Zr1Nwf-OWXEXe-UbuQg{margin-left:8px;margin-right:-7px}[dir=rtl] .jR8x9d .Vo0FCd .VfPpkd-Zr1Nwf-OWXEXe-UbuQg,.jR8x9d .Vo0FCd .VfPpkd-Zr1Nwf-OWXEXe-UbuQg[dir=rtl]{margin-left:-7px;margin-right:8px}.jR8x9d .Vo0FCd .VfPpkd-v1cqY{top:-1px;left:-1px;border:1px solid transparent}.jR8x9d .Vo0FCd.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd{padding-right:11px;padding-left:11px;border-width:1px;border-color:transparent;border-color:var(--gm-chip-outline-color,transparent)}.jR8x9d .Vo0FCd.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd:focus,.jR8x9d .Vo0FCd.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd.VfPpkd-XPtOyb-OWXEXe-ssJRIf-JIbuQc-XpnDCe{padding-right:11px;padding-left:11px;border-width:1px}.jR8x9d .Vo0FCd.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd:focus .VfPpkd-v1cqY,.jR8x9d .Vo0FCd.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd.VfPpkd-XPtOyb-OWXEXe-ssJRIf-JIbuQc-XpnDCe .VfPpkd-v1cqY{top:-1px;left:-1px;border:1px solid transparent}.jR8x9d .Vo0FCd.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-v1cqY{top:-1px;left:-1px;border:1px solid transparent}.jR8x9d .Vo0FCd.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd:focus,.jR8x9d .Vo0FCd.ALA4kc.VfPpkd-XPtOyb-OWXEXe-gk6SMd.VfPpkd-XPtOyb-OWXEXe-ssJRIf-JIbuQc-XpnDCe{border-color:transparent;border-color:var(--gm-chip-outline-color--stateful,transparent)}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-to915-Ia7Qfc .VfPpkd-rOvkhd-Zr1Nwf-OWXEXe-ssJRIf{color:rgb(154,160,166)}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-to915-Ia7Qfc .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf:not(.VfPpkd-rOvkhd-jPmIDe-OWXEXe-SdanKc):hover .VfPpkd-rOvkhd-Zr1Nwf-OWXEXe-ssJRIf{color:rgb(232,234,237)}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-to915-Ia7Qfc .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf:not(.VfPpkd-rOvkhd-jPmIDe-OWXEXe-SdanKc).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-rOvkhd-Zr1Nwf-OWXEXe-ssJRIf,.jR8x9d .UMrnmb-XPtOyb-OWXEXe-to915-Ia7Qfc .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf:not(.VfPpkd-rOvkhd-jPmIDe-OWXEXe-SdanKc):not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-rOvkhd-Zr1Nwf-OWXEXe-ssJRIf{color:rgb(232,234,237)}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-to915-Ia7Qfc.VfPpkd-rOvkhd-XPtOyb-OWXEXe-OWB6Me .VfPpkd-rOvkhd-Zr1Nwf-OWXEXe-ssJRIf{color:rgba(232,234,237,.38)}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-to915-Ia7Qfc .VfPpkd-rOvkhd-TfeOUb-V67aGc{color:rgb(154,160,166)}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-to915-Ia7Qfc .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf:not(.VfPpkd-rOvkhd-jPmIDe-OWXEXe-SdanKc):hover .VfPpkd-rOvkhd-TfeOUb-V67aGc{color:rgb(232,234,237)}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-to915-Ia7Qfc .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf:not(.VfPpkd-rOvkhd-jPmIDe-OWXEXe-SdanKc).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-rOvkhd-TfeOUb-V67aGc,.jR8x9d .UMrnmb-XPtOyb-OWXEXe-to915-Ia7Qfc .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf:not(.VfPpkd-rOvkhd-jPmIDe-OWXEXe-SdanKc):not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-rOvkhd-TfeOUb-V67aGc{color:rgb(232,234,237)}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-to915-Ia7Qfc.VfPpkd-rOvkhd-XPtOyb-OWXEXe-OWB6Me .VfPpkd-rOvkhd-TfeOUb-V67aGc{color:rgba(232,234,237,.38)}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-to915-Ia7Qfc .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf .VfPpkd-rOvkhd-v1cqY::before,.jR8x9d .UMrnmb-XPtOyb-OWXEXe-to915-Ia7Qfc .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf .VfPpkd-rOvkhd-v1cqY::after{background-color:rgb(232,234,237);background-color:var(--mdc-ripple-color,rgb(232,234,237))}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-to915-Ia7Qfc .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf:hover .VfPpkd-rOvkhd-v1cqY::before,.jR8x9d .UMrnmb-XPtOyb-OWXEXe-to915-Ia7Qfc .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-rOvkhd-v1cqY::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-to915-Ia7Qfc .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-rOvkhd-v1cqY::before,.jR8x9d .UMrnmb-XPtOyb-OWXEXe-to915-Ia7Qfc .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-rOvkhd-v1cqY::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-to915-Ia7Qfc .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-rOvkhd-v1cqY::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-to915-Ia7Qfc .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-rOvkhd-v1cqY::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-to915-Ia7Qfc .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-OmTp3c-to915-Ia7Qfc .VfPpkd-rOvkhd-Zr1Nwf-OWXEXe-ssJRIf{color:rgb(138,180,248)}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-OmTp3c-to915-Ia7Qfc .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf:not(.VfPpkd-rOvkhd-jPmIDe-OWXEXe-SdanKc):hover .VfPpkd-rOvkhd-Zr1Nwf-OWXEXe-ssJRIf{color:rgb(138,180,248)}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-OmTp3c-to915-Ia7Qfc .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf:not(.VfPpkd-rOvkhd-jPmIDe-OWXEXe-SdanKc).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-rOvkhd-Zr1Nwf-OWXEXe-ssJRIf,.jR8x9d .UMrnmb-XPtOyb-OWXEXe-OmTp3c-to915-Ia7Qfc .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf:not(.VfPpkd-rOvkhd-jPmIDe-OWXEXe-SdanKc):not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-rOvkhd-Zr1Nwf-OWXEXe-ssJRIf{color:rgb(138,180,248)}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-OmTp3c-to915-Ia7Qfc.VfPpkd-rOvkhd-XPtOyb-OWXEXe-OWB6Me .VfPpkd-rOvkhd-Zr1Nwf-OWXEXe-ssJRIf{color:rgba(232,234,237,.38)}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-OmTp3c-to915-Ia7Qfc .VfPpkd-rOvkhd-TfeOUb-V67aGc{color:rgb(232,234,237)}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-yOOK0-to915-Ia7Qfc.VfPpkd-rOvkhd-XPtOyb-OWXEXe-gk6SMd{background-color:rgba(138,180,248,.24)}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-yOOK0-to915-Ia7Qfc.VfPpkd-rOvkhd-XPtOyb-OWXEXe-gk6SMd.VfPpkd-rOvkhd-XPtOyb-OWXEXe-OWB6Me{background-color:rgba(232,234,237,.12)}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-yOOK0-to915-Ia7Qfc.VfPpkd-rOvkhd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf:before{border-color:transparent}}@media screen and (prefers-color-scheme:dark) and (forced-colors:active){.jR8x9d .UMrnmb-XPtOyb-OWXEXe-yOOK0-to915-Ia7Qfc.VfPpkd-rOvkhd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf:before{border-color:CanvasText}}@media screen and (prefers-color-scheme:dark){.jR8x9d .UMrnmb-XPtOyb-OWXEXe-yOOK0-to915-Ia7Qfc.VfPpkd-rOvkhd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf:not(.VfPpkd-rOvkhd-jPmIDe-OWXEXe-SdanKc).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:before,.jR8x9d .UMrnmb-XPtOyb-OWXEXe-yOOK0-to915-Ia7Qfc.VfPpkd-rOvkhd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf:not(.VfPpkd-rOvkhd-jPmIDe-OWXEXe-SdanKc):not(.VfPpkd-ksKsZd-mWPk3d):focus:before{border-color:transparent}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-yOOK0-to915-Ia7Qfc.VfPpkd-rOvkhd-XPtOyb-OWXEXe-gk6SMd.VfPpkd-rOvkhd-XPtOyb-OWXEXe-OWB6Me .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf:before{border-color:transparent}}@media screen and (prefers-color-scheme:dark) and (forced-colors:active){.jR8x9d .UMrnmb-XPtOyb-OWXEXe-yOOK0-to915-Ia7Qfc.VfPpkd-rOvkhd-XPtOyb-OWXEXe-gk6SMd.VfPpkd-rOvkhd-XPtOyb-OWXEXe-OWB6Me .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf:before{border-color:CanvasText}}@media screen and (prefers-color-scheme:dark){.jR8x9d .UMrnmb-XPtOyb-OWXEXe-yOOK0-to915-Ia7Qfc.VfPpkd-rOvkhd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-rOvkhd-TfeOUb-V67aGc{color:rgb(210,227,252)}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-yOOK0-to915-Ia7Qfc.VfPpkd-rOvkhd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf:not(.VfPpkd-rOvkhd-jPmIDe-OWXEXe-SdanKc):hover .VfPpkd-rOvkhd-TfeOUb-V67aGc{color:#fff}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-yOOK0-to915-Ia7Qfc.VfPpkd-rOvkhd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf:not(.VfPpkd-rOvkhd-jPmIDe-OWXEXe-SdanKc).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-rOvkhd-TfeOUb-V67aGc,.jR8x9d .UMrnmb-XPtOyb-OWXEXe-yOOK0-to915-Ia7Qfc.VfPpkd-rOvkhd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf:not(.VfPpkd-rOvkhd-jPmIDe-OWXEXe-SdanKc):not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-rOvkhd-TfeOUb-V67aGc{color:#fff}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-yOOK0-to915-Ia7Qfc.VfPpkd-rOvkhd-XPtOyb-OWXEXe-gk6SMd.VfPpkd-rOvkhd-XPtOyb-OWXEXe-OWB6Me .VfPpkd-rOvkhd-TfeOUb-V67aGc{color:rgba(232,234,237,.38)}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-yOOK0-to915-Ia7Qfc .VfPpkd-rOvkhd-PvL5qd{color:rgb(210,227,252)}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-yOOK0-to915-Ia7Qfc .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf:not(.VfPpkd-rOvkhd-jPmIDe-OWXEXe-SdanKc):hover .VfPpkd-rOvkhd-PvL5qd{color:#fff}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-yOOK0-to915-Ia7Qfc .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-rOvkhd-PvL5qd,.jR8x9d .UMrnmb-XPtOyb-OWXEXe-yOOK0-to915-Ia7Qfc .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-rOvkhd-PvL5qd{color:#fff}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-yOOK0-to915-Ia7Qfc.VfPpkd-rOvkhd-XPtOyb-OWXEXe-OWB6Me .VfPpkd-rOvkhd-PvL5qd{color:rgba(232,234,237,.38)}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-yOOK0-to915-Ia7Qfc.VfPpkd-rOvkhd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf .VfPpkd-rOvkhd-v1cqY::before,.jR8x9d .UMrnmb-XPtOyb-OWXEXe-yOOK0-to915-Ia7Qfc.VfPpkd-rOvkhd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf .VfPpkd-rOvkhd-v1cqY::after{background-color:#fff;background-color:var(--mdc-ripple-color,#fff)}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-yOOK0-to915-Ia7Qfc.VfPpkd-rOvkhd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf:hover .VfPpkd-rOvkhd-v1cqY::before,.jR8x9d .UMrnmb-XPtOyb-OWXEXe-yOOK0-to915-Ia7Qfc.VfPpkd-rOvkhd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-rOvkhd-v1cqY::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-yOOK0-to915-Ia7Qfc.VfPpkd-rOvkhd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-rOvkhd-v1cqY::before,.jR8x9d .UMrnmb-XPtOyb-OWXEXe-yOOK0-to915-Ia7Qfc.VfPpkd-rOvkhd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-rOvkhd-v1cqY::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-yOOK0-to915-Ia7Qfc.VfPpkd-rOvkhd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-rOvkhd-v1cqY::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-yOOK0-to915-Ia7Qfc.VfPpkd-rOvkhd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-rOvkhd-v1cqY::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-yOOK0-to915-Ia7Qfc.VfPpkd-rOvkhd-XPtOyb-OWXEXe-gk6SMd .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-YPqjbf-to915-Ia7Qfc .VfPpkd-rOvkhd-Zr1Nwf-OWXEXe-UbuQg{color:rgb(154,160,166)}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-YPqjbf-to915-Ia7Qfc .VfPpkd-rOvkhd-jPmIDe-OWXEXe-UbuQg:hover .VfPpkd-rOvkhd-Zr1Nwf-OWXEXe-UbuQg{color:rgb(232,234,237)}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-YPqjbf-to915-Ia7Qfc .VfPpkd-rOvkhd-jPmIDe-OWXEXe-UbuQg.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-rOvkhd-Zr1Nwf-OWXEXe-UbuQg,.jR8x9d .UMrnmb-XPtOyb-OWXEXe-YPqjbf-to915-Ia7Qfc .VfPpkd-rOvkhd-jPmIDe-OWXEXe-UbuQg:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-rOvkhd-Zr1Nwf-OWXEXe-UbuQg{color:rgb(232,234,237)}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-YPqjbf-to915-Ia7Qfc.VfPpkd-rOvkhd-XPtOyb-OWXEXe-OWB6Me .VfPpkd-rOvkhd-Zr1Nwf-OWXEXe-UbuQg{color:rgba(232,234,237,.38)}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-YPqjbf-to915-Ia7Qfc .VfPpkd-rOvkhd-jPmIDe-OWXEXe-UbuQg .VfPpkd-rOvkhd-v1cqY::before,.jR8x9d .UMrnmb-XPtOyb-OWXEXe-YPqjbf-to915-Ia7Qfc .VfPpkd-rOvkhd-jPmIDe-OWXEXe-UbuQg .VfPpkd-rOvkhd-v1cqY::after{background-color:rgb(232,234,237);background-color:var(--mdc-ripple-color,rgb(232,234,237))}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-YPqjbf-to915-Ia7Qfc .VfPpkd-rOvkhd-jPmIDe-OWXEXe-UbuQg:hover .VfPpkd-rOvkhd-v1cqY::before,.jR8x9d .UMrnmb-XPtOyb-OWXEXe-YPqjbf-to915-Ia7Qfc .VfPpkd-rOvkhd-jPmIDe-OWXEXe-UbuQg.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-rOvkhd-v1cqY::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-YPqjbf-to915-Ia7Qfc .VfPpkd-rOvkhd-jPmIDe-OWXEXe-UbuQg.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-rOvkhd-v1cqY::before,.jR8x9d .UMrnmb-XPtOyb-OWXEXe-YPqjbf-to915-Ia7Qfc .VfPpkd-rOvkhd-jPmIDe-OWXEXe-UbuQg:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-rOvkhd-v1cqY::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-YPqjbf-to915-Ia7Qfc .VfPpkd-rOvkhd-jPmIDe-OWXEXe-UbuQg:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-rOvkhd-v1cqY::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-YPqjbf-to915-Ia7Qfc .VfPpkd-rOvkhd-jPmIDe-OWXEXe-UbuQg:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-rOvkhd-v1cqY::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-YPqjbf-to915-Ia7Qfc .VfPpkd-rOvkhd-jPmIDe-OWXEXe-UbuQg.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-aSvl1d-to915-Ia7Qfc{background-color:transparent}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-aSvl1d-to915-Ia7Qfc .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf:before{border-width:1px}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-aSvl1d-to915-Ia7Qfc .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf:before{border-style:solid}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-aSvl1d-to915-Ia7Qfc.VfPpkd-rOvkhd-XPtOyb-OWXEXe-OWB6Me{background-color:transparent}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-aSvl1d-to915-Ia7Qfc .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf:before{border-color:rgb(95,99,104)}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-aSvl1d-to915-Ia7Qfc .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf:not(.VfPpkd-rOvkhd-jPmIDe-OWXEXe-SdanKc).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:before,.jR8x9d .UMrnmb-XPtOyb-OWXEXe-aSvl1d-to915-Ia7Qfc .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf:not(.VfPpkd-rOvkhd-jPmIDe-OWXEXe-SdanKc):not(.VfPpkd-ksKsZd-mWPk3d):focus:before{border-color:rgb(232,234,237)}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-aSvl1d-to915-Ia7Qfc.VfPpkd-rOvkhd-XPtOyb-OWXEXe-OWB6Me .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf:before{border-color:rgba(232,234,237,.12)}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-ITYOJe-to915-Ia7Qfc{background-color:rgb(32,33,36);-webkit-transition:border .28s cubic-bezier(.4,0,.2,1),box-shadow .28s cubic-bezier(.4,0,.2,1);transition:border .28s cubic-bezier(.4,0,.2,1),box-shadow .28s cubic-bezier(.4,0,.2,1);box-shadow:0 1px 2px 0 rgba(0,0,0,.3),0 1px 3px 1px rgba(0,0,0,.15)}}@media screen and (prefers-color-scheme:dark) and (-ms-high-contrast:active),screen and (prefers-color-scheme:dark) and (forced-colors:active){.jR8x9d .UMrnmb-XPtOyb-OWXEXe-ITYOJe-to915-Ia7Qfc .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf:before{border-width:1px}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-ITYOJe-to915-Ia7Qfc .VfPpkd-rOvkhd-jPmIDe-OWXEXe-ssJRIf:before{border-style:solid}}@media screen and (prefers-color-scheme:dark){.jR8x9d .UMrnmb-XPtOyb-OWXEXe-ITYOJe-to915-Ia7Qfc.VfPpkd-rOvkhd-XPtOyb-OWXEXe-OWB6Me{background-color:rgba(232,234,237,.12)}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-ITYOJe-to915-Ia7Qfc .VfPpkd-BFbNVe-bF1uUb{opacity:.05}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-ITYOJe-to915-Ia7Qfc:hover{box-shadow:0 1px 2px 0 rgba(0,0,0,.3),0 2px 6px 2px rgba(0,0,0,.15)}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-ITYOJe-to915-Ia7Qfc:hover .VfPpkd-BFbNVe-bF1uUb{opacity:.08}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-ITYOJe-to915-Ia7Qfc:active{box-shadow:0 1px 3px 0 rgba(0,0,0,.3),0 4px 8px 3px rgba(0,0,0,.15)}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-ITYOJe-to915-Ia7Qfc:active .VfPpkd-BFbNVe-bF1uUb{opacity:.11}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-ITYOJe-to915-Ia7Qfc.VfPpkd-rOvkhd-XPtOyb-OWXEXe-OWB6Me{box-shadow:none}.jR8x9d .UMrnmb-XPtOyb-OWXEXe-ITYOJe-to915-Ia7Qfc.VfPpkd-rOvkhd-XPtOyb-OWXEXe-OWB6Me .VfPpkd-BFbNVe-bF1uUb{opacity:0}.jR8x9d .a9u1Hb .VfPpkd-JGcpL-uI4vCe-LkdAo,.jR8x9d .a9u1Hb .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:rgb(102,157,246)}}@media screen and (prefers-color-scheme:dark) and (-ms-high-contrast:active),screen and (prefers-color-scheme:dark) and (forced-colors:active){.jR8x9d .a9u1Hb .VfPpkd-JGcpL-uI4vCe-LkdAo,.jR8x9d .a9u1Hb .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:CanvasText}}@media screen and (prefers-color-scheme:dark){.jR8x9d .a9u1Hb .VfPpkd-JGcpL-Ydhldb-R6PoUb .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:rgb(66,133,244)}}@media screen and (prefers-color-scheme:dark) and (-ms-high-contrast:active),screen and (prefers-color-scheme:dark) and (forced-colors:active){.jR8x9d .a9u1Hb .VfPpkd-JGcpL-Ydhldb-R6PoUb .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:CanvasText}}@media screen and (prefers-color-scheme:dark){.jR8x9d .a9u1Hb .VfPpkd-JGcpL-Ydhldb-ibL1re .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:rgb(234,67,53)}}@media screen and (prefers-color-scheme:dark) and (-ms-high-contrast:active),screen and (prefers-color-scheme:dark) and (forced-colors:active){.jR8x9d .a9u1Hb .VfPpkd-JGcpL-Ydhldb-ibL1re .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:CanvasText}}@media screen and (prefers-color-scheme:dark){.jR8x9d .a9u1Hb .VfPpkd-JGcpL-Ydhldb-c5RTEf .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:rgb(251,188,4)}}@media screen and (prefers-color-scheme:dark) and (-ms-high-contrast:active),screen and (prefers-color-scheme:dark) and (forced-colors:active){.jR8x9d .a9u1Hb .VfPpkd-JGcpL-Ydhldb-c5RTEf .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:CanvasText}}@media screen and (prefers-color-scheme:dark){.jR8x9d .a9u1Hb .VfPpkd-JGcpL-Ydhldb-II5mzb .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:rgb(52,168,83)}}@media screen and (prefers-color-scheme:dark) and (-ms-high-contrast:active),screen and (prefers-color-scheme:dark) and (forced-colors:active){.jR8x9d .a9u1Hb .VfPpkd-JGcpL-Ydhldb-II5mzb .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:CanvasText}}@media screen and (prefers-color-scheme:dark){.jR8x9d .tKSZFd{background-color:rgb(32,33,36);border-color:rgb(95,99,104)}.jR8x9d .tKSZFd .VfPpkd-wZVHld-vqLbZd-eEDwDf{background-color:rgb(32,33,36)}.jR8x9d .tKSZFd .VfPpkd-wZVHld-vqLbZd-eEDwDf,.jR8x9d .tKSZFd .VfPpkd-wZVHld-gruSEe-j4LONd,.jR8x9d .tKSZFd .VfPpkd-wZVHld-gruSEe-YMi5E-I8r9Db-DARUcf-V67aGc,.jR8x9d .tKSZFd .VfPpkd-wZVHld-aOtOmf{color:rgb(232,234,237)}.jR8x9d .tKSZFd .VfPpkd-wZVHld-xMbwt-OWXEXe-gk6SMd{background-color:rgba(138,180,248,.24)}.jR8x9d .tKSZFd .VfPpkd-wZVHld-gruSEe-YMi5E-I8r9Db-DARUcf-O1htCb-OWXEXe-INsAgc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Brv4Fb,.jR8x9d .tKSZFd .VfPpkd-wZVHld-gruSEe-YMi5E-I8r9Db-DARUcf-O1htCb-OWXEXe-INsAgc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Ra9xwd,.jR8x9d .tKSZFd .VfPpkd-wZVHld-gruSEe-YMi5E-I8r9Db-DARUcf-O1htCb-OWXEXe-INsAgc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-MpmGFe{border-color:rgb(95,99,104)}.jR8x9d .tKSZFd .VfPpkd-wZVHld-aOtOmf,.jR8x9d .tKSZFd .VfPpkd-wZVHld-vqLbZd-eEDwDf{border-bottom-color:rgb(95,99,104)}.jR8x9d .tKSZFd .VfPpkd-wZVHld-gruSEe{border-top-color:rgb(95,99,104)}.jR8x9d .tKSZFd .VfPpkd-wZVHld-xMbwt:not(.VfPpkd-wZVHld-xMbwt-OWXEXe-gk6SMd):hover{background-color:rgba(232,234,237,.04)}.jR8x9d .tKSZFd .VfPpkd-wZVHld-EcJZQc-Bz112c-LgbsSe{color:rgb(154,160,166)}.jR8x9d .tKSZFd .VfPpkd-wZVHld-EcJZQc-Bz112c-LgbsSe .VfPpkd-Bz112c-Jh9lGc::before,.jR8x9d .tKSZFd .VfPpkd-wZVHld-EcJZQc-Bz112c-LgbsSe .VfPpkd-Bz112c-Jh9lGc::after{background-color:rgb(154,160,166);background-color:var(--mdc-ripple-color,rgb(154,160,166))}.jR8x9d .tKSZFd .VfPpkd-wZVHld-EcJZQc-Bz112c-LgbsSe:hover .VfPpkd-Bz112c-Jh9lGc::before,.jR8x9d .tKSZFd .VfPpkd-wZVHld-EcJZQc-Bz112c-LgbsSe.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Bz112c-Jh9lGc::before{opacity:.08;opacity:var(--mdc-ripple-hover-opacity,.08)}.jR8x9d .tKSZFd .VfPpkd-wZVHld-EcJZQc-Bz112c-LgbsSe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Bz112c-Jh9lGc::before,.jR8x9d .tKSZFd .VfPpkd-wZVHld-EcJZQc-Bz112c-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Bz112c-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.24;opacity:var(--mdc-ripple-focus-opacity,.24)}.jR8x9d .tKSZFd .VfPpkd-wZVHld-EcJZQc-Bz112c-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Bz112c-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .tKSZFd .VfPpkd-wZVHld-EcJZQc-Bz112c-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Bz112c-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.24;opacity:var(--mdc-ripple-press-opacity,.24)}.jR8x9d .tKSZFd .VfPpkd-wZVHld-EcJZQc-Bz112c-LgbsSe.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.24)}.jR8x9d .tKSZFd .VfPpkd-wZVHld-vqLbZd-eEDwDf-OWXEXe-Evexob .VfPpkd-wZVHld-EcJZQc-Bz112c-LgbsSe{color:rgb(232,234,237)}.jR8x9d .tKSZFd .VfPpkd-wZVHld-vqLbZd-eEDwDf-OWXEXe-Evexob .VfPpkd-wZVHld-EcJZQc-Bz112c-LgbsSe .VfPpkd-Bz112c-Jh9lGc::before,.jR8x9d .tKSZFd .VfPpkd-wZVHld-vqLbZd-eEDwDf-OWXEXe-Evexob .VfPpkd-wZVHld-EcJZQc-Bz112c-LgbsSe .VfPpkd-Bz112c-Jh9lGc::after{background-color:rgb(232,234,237);background-color:var(--mdc-ripple-color,rgb(232,234,237))}.jR8x9d .tKSZFd .VfPpkd-wZVHld-vqLbZd-eEDwDf-OWXEXe-Evexob .VfPpkd-wZVHld-EcJZQc-Bz112c-LgbsSe:hover .VfPpkd-Bz112c-Jh9lGc::before,.jR8x9d .tKSZFd .VfPpkd-wZVHld-vqLbZd-eEDwDf-OWXEXe-Evexob .VfPpkd-wZVHld-EcJZQc-Bz112c-LgbsSe.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Bz112c-Jh9lGc::before{opacity:.08;opacity:var(--mdc-ripple-hover-opacity,.08)}.jR8x9d .tKSZFd .VfPpkd-wZVHld-vqLbZd-eEDwDf-OWXEXe-Evexob .VfPpkd-wZVHld-EcJZQc-Bz112c-LgbsSe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Bz112c-Jh9lGc::before,.jR8x9d .tKSZFd .VfPpkd-wZVHld-vqLbZd-eEDwDf-OWXEXe-Evexob .VfPpkd-wZVHld-EcJZQc-Bz112c-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Bz112c-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.24;opacity:var(--mdc-ripple-focus-opacity,.24)}.jR8x9d .tKSZFd .VfPpkd-wZVHld-vqLbZd-eEDwDf-OWXEXe-Evexob .VfPpkd-wZVHld-EcJZQc-Bz112c-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Bz112c-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .tKSZFd .VfPpkd-wZVHld-vqLbZd-eEDwDf-OWXEXe-Evexob .VfPpkd-wZVHld-EcJZQc-Bz112c-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Bz112c-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.24;opacity:var(--mdc-ripple-press-opacity,.24)}.jR8x9d .tKSZFd .VfPpkd-wZVHld-vqLbZd-eEDwDf-OWXEXe-Evexob .VfPpkd-wZVHld-EcJZQc-Bz112c-LgbsSe.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.24)}.jR8x9d .zNgRPc .bwNLcf{color:rgb(232,234,237);font-family:Roboto,Arial,sans-serif;line-height:1.5rem;font-size:1rem;letter-spacing:.00625em;font-weight:400}.jR8x9d .zNgRPc .bwNLcf .VfPpkd-StrnGf-rymPhb-IhFlZd{color:rgb(154,160,166)}.jR8x9d .zNgRPc .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS{color:rgb(232,234,237)}.jR8x9d .zNgRPc .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c{opacity:.38}.jR8x9d .zNgRPc .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-f7MjDc,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-f7MjDc{color:rgb(232,234,237)}.jR8x9d .zNgRPc .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:0}.jR8x9d .zNgRPc .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd{background-color:rgba(138,180,248,.24)}.jR8x9d .zNgRPc .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::after{background-color:rgb(138,180,248);background-color:var(--mdc-ripple-color,rgb(138,180,248))}.jR8x9d .zNgRPc .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.jR8x9d .zNgRPc .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.jR8x9d .zNgRPc .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .zNgRPc .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.jR8x9d .zNgRPc .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}.jR8x9d .zNgRPc .bwNLcf .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS{color:rgb(154,160,166)}.jR8x9d .zNgRPc .bwNLcf .VfPpkd-StrnGf-rymPhb-clz4Ic{border-bottom-color:rgba(232,234,237,.12)}.jR8x9d .zNgRPc .bwNLcf .VfPpkd-StrnGf-rymPhb-f7MjDc{color:rgb(232,234,237)}.jR8x9d .zNgRPc .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-pZXsl::before,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-pZXsl::after{background-color:rgb(232,234,237);background-color:var(--mdc-ripple-color,rgb(232,234,237))}.jR8x9d .zNgRPc .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.jR8x9d .zNgRPc .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.jR8x9d .zNgRPc .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .zNgRPc .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.jR8x9d .zNgRPc .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}}@media screen and (prefers-color-scheme:dark) and (-ms-high-contrast:active),screen and (prefers-color-scheme:dark) and (forced-colors:active){.jR8x9d .zNgRPc .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS{color:GrayText}.jR8x9d .zNgRPc .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c{opacity:1}}@media screen and (prefers-color-scheme:dark){.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-Gtdoyb,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-fpDzbe-fmcmS{color:rgb(232,234,237)}.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-L8ivfd-fmcmS,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-bC5pod-fmcmS,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-JMEf7e{color:rgb(154,160,166)}.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-Gtdoyb,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-fpDzbe-fmcmS,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-L8ivfd-fmcmS,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-bC5pod-fmcmS,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e{color:rgb(232,234,237)}.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-KkROqb,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-Gtdoyb,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-JMEf7e{opacity:.38}.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-Gtdoyb,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-fpDzbe-fmcmS,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-rymPhb-Gtdoyb,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-rymPhb-fpDzbe-fmcmS,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb{color:rgb(232,234,237)}.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::before{opacity:0}.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd{background-color:rgba(138,180,248,.24)}.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::before,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::after{background-color:rgb(138,180,248);background-color:var(--mdc-ripple-color,rgb(138,180,248))}.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-rymPhb-pZXsl::before,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-rymPhb-pZXsl::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-rymPhb-pZXsl::before,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-rymPhb-pZXsl::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-rymPhb-pZXsl::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-rymPhb-pZXsl::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-L8ivfd-fmcmS{color:rgb(154,160,166)}.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-clz4Ic{background-color:rgba(232,234,237,.12)}.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e{color:rgb(232,234,237)}.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::before,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::after{background-color:rgb(232,234,237);background-color:var(--mdc-ripple-color,rgb(232,234,237))}.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b:hover .VfPpkd-rymPhb-pZXsl::before,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-rymPhb-pZXsl::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-rymPhb-pZXsl::before,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-rymPhb-pZXsl::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-rymPhb-pZXsl::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-rymPhb-pZXsl::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}}@media screen and (prefers-color-scheme:dark) and (forced-colors:active){.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-Gtdoyb,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-fpDzbe-fmcmS,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-L8ivfd-fmcmS,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-bC5pod-fmcmS,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e{color:GrayText}.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-KkROqb,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-Gtdoyb,.jR8x9d .zNgRPc .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-JMEf7e{opacity:1}}@media screen and (prefers-color-scheme:dark){.jR8x9d .zNgRPc .VfPpkd-XqMb-hFsbo{color:rgb(154,160,166)}.jR8x9d .zNgRPc .VfPpkd-XqMb-hFsbo:hover{color:rgb(248,249,250)}.jR8x9d .zNgRPc .VfPpkd-XqMb-hFsbo.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.jR8x9d .zNgRPc .VfPpkd-XqMb-hFsbo:not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(248,249,250)}.jR8x9d .zNgRPc .VfPpkd-XqMb-hFsbo:not(:disabled):active{color:rgb(248,249,250)}.jR8x9d .zNgRPc .VfPpkd-XqMb-hFsbo .VfPpkd-Bz112c-Jh9lGc::before,.jR8x9d .zNgRPc .VfPpkd-XqMb-hFsbo .VfPpkd-Bz112c-Jh9lGc::after{background-color:rgb(232,234,237);background-color:var(--mdc-ripple-color,rgb(232,234,237))}.jR8x9d .zNgRPc .VfPpkd-XqMb-hFsbo-OWXEXe-FGU2Pb-OWB6Me{color:rgba(232,234,237,.38)}.jR8x9d .zNgRPc .VfPpkd-XqMb-hFsbo-OWXEXe-FGU2Pb-OWB6Me:hover,.jR8x9d .zNgRPc .VfPpkd-XqMb-hFsbo-OWXEXe-FGU2Pb-OWB6Me.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.jR8x9d .zNgRPc .VfPpkd-XqMb-hFsbo-OWXEXe-FGU2Pb-OWB6Me:not(.VfPpkd-ksKsZd-mWPk3d):focus,.jR8x9d .zNgRPc .VfPpkd-XqMb-hFsbo-OWXEXe-FGU2Pb-OWB6Me:not(:disabled):active{color:rgba(232,234,237,.38)}.jR8x9d .zNgRPc .VfPpkd-XqMb-S2QgGf-kj0dLd:not(:disabled){color:rgb(154,160,166);color:var(--mdc-text-button-label-text-color,rgb(154,160,166))}.jR8x9d .zNgRPc .VfPpkd-XqMb-S2QgGf-kj0dLd:not(:disabled):hover{color:rgb(248,249,250);color:var(--mdc-text-button-hover-label-text-color,rgb(248,249,250))}.jR8x9d .zNgRPc .VfPpkd-XqMb-S2QgGf-kj0dLd:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.jR8x9d .zNgRPc .VfPpkd-XqMb-S2QgGf-kj0dLd:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(248,249,250);color:var(--mdc-text-button-focus-label-text-color,rgb(248,249,250))}.jR8x9d .zNgRPc .VfPpkd-XqMb-S2QgGf-kj0dLd:not(:disabled):not(:disabled):active{color:rgb(248,249,250);color:var(--mdc-text-button-pressed-label-text-color,rgb(248,249,250))}.jR8x9d .zNgRPc .VfPpkd-XqMb-S2QgGf-kj0dLd:disabled{color:rgb(154,160,166);color:var(--mdc-text-button-disabled-label-text-color,rgb(154,160,166))}.jR8x9d .zNgRPc .VfPpkd-hOoMI-haAclf .VfPpkd-hOoMI-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd{background-color:transparent}.jR8x9d .zNgRPc .VfPpkd-hOoMI-haAclf .VfPpkd-hOoMI-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::before,.jR8x9d .zNgRPc .VfPpkd-hOoMI-haAclf .VfPpkd-hOoMI-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::after{background-color:rgb(232,234,237);background-color:var(--mdc-ripple-color,rgb(232,234,237))}.jR8x9d .zNgRPc .VfPpkd-hOoMI-haAclf{background-color:rgb(32,33,36)}.jR8x9d .zNgRPc.VfPpkd-Zc28rc-OWXEXe-Mgvhmd-S2QgGf-FNFY6c .VfPpkd-XqMb-S2QgGf-kj0dLd:not(:disabled),.jR8x9d .zNgRPc.VfPpkd-Zc28rc-OWXEXe-WRCQcd-S2QgGf-FNFY6c .VfPpkd-XqMb-S2QgGf-kj0dLd:not(:disabled){color:rgb(248,249,250);color:var(--mdc-text-button-label-text-color,rgb(248,249,250))}.jR8x9d .zNgRPc.VfPpkd-Zc28rc-OWXEXe-Mgvhmd-S2QgGf-FNFY6c .VfPpkd-XqMb-S2QgGf-kj0dLd:not(:disabled),.jR8x9d .zNgRPc.VfPpkd-Zc28rc-OWXEXe-WRCQcd-S2QgGf-FNFY6c .VfPpkd-XqMb-S2QgGf-kj0dLd:not(:disabled){background-color:rgba(232,234,237,.12)}.jR8x9d .zNgRPc.VfPpkd-Zc28rc-OWXEXe-Mgvhmd-S2QgGf-FNFY6c .VfPpkd-hOoMI-haAclf,.jR8x9d .zNgRPc.VfPpkd-Zc28rc-OWXEXe-WRCQcd-S2QgGf-FNFY6c .VfPpkd-hOoMI-haAclf{border-top-color:rgb(95,99,104)}.jR8x9d .zNgRPc .VfPpkd-HhDot-tJHJj{color:rgb(154,160,166)}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe:not(:disabled){color:rgb(232,234,237);color:var(--mdc-outlined-button-label-text-color,rgb(232,234,237))}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe:not(:disabled):hover{color:rgb(248,249,250);color:var(--mdc-outlined-button-hover-label-text-color,rgb(248,249,250))}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(248,249,250);color:var(--mdc-outlined-button-focus-label-text-color,rgb(248,249,250))}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe:not(:disabled):not(:disabled):active{color:rgb(248,249,250);color:var(--mdc-outlined-button-pressed-label-text-color,rgb(248,249,250))}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe:disabled{color:rgb(154,160,166);color:var(--mdc-outlined-button-disabled-label-text-color,rgb(154,160,166))}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe .VfPpkd-Jh9lGc::before{background-color:rgb(232,234,237);background-color:var(--mdc-outlined-button-hover-state-layer-color,rgb(232,234,237))}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe .VfPpkd-Jh9lGc::after{background-color:rgb(232,234,237);background-color:var(--mdc-outlined-button-pressed-state-layer-color,rgb(232,234,237))}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe:hover .VfPpkd-Jh9lGc::before,.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:.04;opacity:var(--mdc-outlined-button-hover-state-layer-opacity,.04)}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-outlined-button-focus-state-layer-opacity,.12)}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-outlined-button-pressed-state-layer-opacity,.1)}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-outlined-button-pressed-state-layer-opacity,0.1)}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled){color:rgb(138,180,248);color:var(--mdc-outlined-button-label-text-color,rgb(138,180,248))}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled):hover{color:rgb(174,203,250);color:var(--mdc-outlined-button-hover-label-text-color,rgb(174,203,250))}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(174,203,250);color:var(--mdc-outlined-button-focus-label-text-color,rgb(174,203,250))}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled):not(:disabled):active{color:rgb(174,203,250);color:var(--mdc-outlined-button-pressed-label-text-color,rgb(174,203,250))}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l .VfPpkd-Jh9lGc::before{background-color:rgb(174,203,250);background-color:var(--mdc-outlined-button-hover-state-layer-color,rgb(174,203,250))}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l .VfPpkd-Jh9lGc::after{background-color:rgb(174,203,250);background-color:var(--mdc-outlined-button-pressed-state-layer-color,rgb(174,203,250))}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:hover .VfPpkd-Jh9lGc::before,.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:.04;opacity:var(--mdc-outlined-button-hover-state-layer-opacity,.04)}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-outlined-button-focus-state-layer-opacity,.12)}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-outlined-button-pressed-state-layer-opacity,.1)}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-outlined-button-pressed-state-layer-opacity,0.1)}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled){border-color:rgb(138,180,248);border-color:var(--mdc-outlined-button-outline-color,rgb(138,180,248))}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{border-color:rgb(174,203,250);border-color:var(--mdc-outlined-button-focus-outline-color,rgb(174,203,250))}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled):hover{border-color:rgb(174,203,250)}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled):active,.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled):focus:active{border-color:rgb(174,203,250)}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(:disabled){color:rgb(32,33,36);color:var(--mdc-outlined-button-label-text-color,rgb(32,33,36))}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(:disabled):hover{color:rgb(32,33,36);color:var(--mdc-outlined-button-hover-label-text-color,rgb(32,33,36))}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(32,33,36);color:var(--mdc-outlined-button-focus-label-text-color,rgb(32,33,36))}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(:disabled):not(:disabled):active{color:rgb(32,33,36);color:var(--mdc-outlined-button-pressed-label-text-color,rgb(32,33,36))}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd .VfPpkd-Jh9lGc::before{background-color:#fff;background-color:var(--mdc-outlined-button-hover-state-layer-color,#fff)}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd .VfPpkd-Jh9lGc::after{background-color:#fff;background-color:var(--mdc-outlined-button-pressed-state-layer-color,#fff)}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:hover .VfPpkd-Jh9lGc::before,.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:.16;opacity:var(--mdc-outlined-button-hover-state-layer-opacity,.16)}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.24;opacity:var(--mdc-outlined-button-focus-state-layer-opacity,.24)}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.2;opacity:var(--mdc-outlined-button-pressed-state-layer-opacity,.2)}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-outlined-button-pressed-state-layer-opacity,0.2)}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(:disabled){background-color:rgb(138,180,248)}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(:disabled):hover{background-color:rgb(138,180,248)}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{background-color:rgb(138,180,248)}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(:disabled):not(:disabled):active{background-color:rgb(138,180,248)}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-OWB6Me:not(:disabled){color:rgb(154,160,166);color:var(--mdc-outlined-button-label-text-color,rgb(154,160,166))}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-OWB6Me:not(:disabled):hover{color:rgb(154,160,166);color:var(--mdc-outlined-button-hover-label-text-color,rgb(154,160,166))}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-OWB6Me:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-OWB6Me:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(154,160,166);color:var(--mdc-outlined-button-focus-label-text-color,rgb(154,160,166))}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-OWB6Me:not(:disabled):not(:disabled):active{color:rgb(154,160,166);color:var(--mdc-outlined-button-pressed-label-text-color,rgb(154,160,166))}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6:not(:disabled){color:rgb(154,160,166);color:var(--mdc-outlined-button-label-text-color,rgb(154,160,166))}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6:not(:disabled):hover{color:rgb(248,249,250);color:var(--mdc-outlined-button-hover-label-text-color,rgb(248,249,250))}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(248,249,250);color:var(--mdc-outlined-button-focus-label-text-color,rgb(248,249,250))}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6:not(:disabled):not(:disabled):active{color:rgb(248,249,250);color:var(--mdc-outlined-button-pressed-label-text-color,rgb(248,249,250))}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled){color:rgb(138,180,248);color:var(--mdc-outlined-button-label-text-color,rgb(138,180,248))}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled):hover{color:rgb(174,203,250);color:var(--mdc-outlined-button-hover-label-text-color,rgb(174,203,250))}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(174,203,250);color:var(--mdc-outlined-button-focus-label-text-color,rgb(174,203,250))}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled):not(:disabled):active{color:rgb(174,203,250);color:var(--mdc-outlined-button-pressed-label-text-color,rgb(174,203,250))}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l .VfPpkd-Jh9lGc::before{background-color:rgb(174,203,250);background-color:var(--mdc-outlined-button-hover-state-layer-color,rgb(174,203,250))}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l .VfPpkd-Jh9lGc::after{background-color:rgb(174,203,250);background-color:var(--mdc-outlined-button-pressed-state-layer-color,rgb(174,203,250))}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:hover .VfPpkd-Jh9lGc::before,.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:.04;opacity:var(--mdc-outlined-button-hover-state-layer-opacity,.04)}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-outlined-button-focus-state-layer-opacity,.12)}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-outlined-button-pressed-state-layer-opacity,.1)}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-outlined-button-pressed-state-layer-opacity,0.1)}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled){border-color:rgb(138,180,248);border-color:var(--mdc-outlined-button-outline-color,rgb(138,180,248))}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{border-color:rgb(174,203,250);border-color:var(--mdc-outlined-button-focus-outline-color,rgb(174,203,250))}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled):hover{border-color:rgb(174,203,250)}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled):active,.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-bAa4l:not(:disabled):focus:active{border-color:rgb(174,203,250)}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(:disabled){color:rgb(32,33,36);color:var(--mdc-outlined-button-label-text-color,rgb(32,33,36))}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(:disabled):hover{color:rgb(32,33,36);color:var(--mdc-outlined-button-hover-label-text-color,rgb(32,33,36))}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(32,33,36);color:var(--mdc-outlined-button-focus-label-text-color,rgb(32,33,36))}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(:disabled):not(:disabled):active{color:rgb(32,33,36);color:var(--mdc-outlined-button-pressed-label-text-color,rgb(32,33,36))}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd .VfPpkd-Jh9lGc::before{background-color:#fff;background-color:var(--mdc-outlined-button-hover-state-layer-color,#fff)}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd .VfPpkd-Jh9lGc::after{background-color:#fff;background-color:var(--mdc-outlined-button-pressed-state-layer-color,#fff)}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:hover .VfPpkd-Jh9lGc::before,.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:.16;opacity:var(--mdc-outlined-button-hover-state-layer-opacity,.16)}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.24;opacity:var(--mdc-outlined-button-focus-state-layer-opacity,.24)}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.2;opacity:var(--mdc-outlined-button-pressed-state-layer-opacity,.2)}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-outlined-button-pressed-state-layer-opacity,0.2)}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(:disabled){background-color:rgb(138,180,248)}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(:disabled):hover{background-color:rgb(138,180,248)}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{background-color:rgb(138,180,248)}.jR8x9d .zNgRPc .VfPpkd-RKhZBe-LgbsSe-OWXEXe-C3kE6.VfPpkd-RKhZBe-LgbsSe-OWXEXe-gk6SMd:not(:disabled):not(:disabled):active{background-color:rgb(138,180,248)}.jR8x9d .f8F5Dd{background-color:rgb(32,33,36);border-width:0;box-shadow:0 1px 2px 0 rgba(0,0,0,.3),0 2px 6px 2px rgba(0,0,0,.15)}.jR8x9d .f8F5Dd .VfPpkd-BFbNVe-bF1uUb{opacity:.08}.jR8x9d .ad0uI .VfPpkd-GRS59e:not(:disabled){color:rgb(138,180,248);color:var(--mdc-text-button-label-text-color,rgb(138,180,248))}.jR8x9d .ad0uI .VfPpkd-GRS59e:not(:disabled):hover{color:rgb(174,203,250);color:var(--mdc-text-button-hover-label-text-color,rgb(174,203,250))}.jR8x9d .ad0uI .VfPpkd-GRS59e:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.jR8x9d .ad0uI .VfPpkd-GRS59e:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(174,203,250);color:var(--mdc-text-button-focus-label-text-color,rgb(174,203,250))}.jR8x9d .ad0uI .VfPpkd-GRS59e:not(:disabled):not(:disabled):active{color:rgb(174,203,250);color:var(--mdc-text-button-pressed-label-text-color,rgb(174,203,250))}.jR8x9d .ad0uI .VfPpkd-GRS59e .VfPpkd-Jh9lGc::before{background-color:rgb(174,203,250);background-color:var(--mdc-text-button-hover-state-layer-color,rgb(174,203,250))}.jR8x9d .ad0uI .VfPpkd-GRS59e .VfPpkd-Jh9lGc::after{background-color:rgb(174,203,250);background-color:var(--mdc-text-button-pressed-state-layer-color,rgb(174,203,250))}.jR8x9d .ad0uI .VfPpkd-GRS59e:hover .VfPpkd-Jh9lGc::before,.jR8x9d .ad0uI .VfPpkd-GRS59e.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:.04;opacity:var(--mdc-text-button-hover-state-layer-opacity,.04)}.jR8x9d .ad0uI .VfPpkd-GRS59e.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.jR8x9d .ad0uI .VfPpkd-GRS59e:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-text-button-focus-state-layer-opacity,.12)}.jR8x9d .ad0uI .VfPpkd-GRS59e:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .ad0uI .VfPpkd-GRS59e:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-text-button-pressed-state-layer-opacity,.1)}.jR8x9d .ad0uI .VfPpkd-GRS59e.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-text-button-pressed-state-layer-opacity,0.1)}.jR8x9d .zF2sRd .VfPpkd-Cv7pCf-ornU0b{color:rgb(189,193,198)}.jR8x9d .zF2sRd .VfPpkd-Cv7pCf-ornU0b:disabled{color:rgba(232,234,237,.38)}.jR8x9d .zF2sRd .VfPpkd-Cv7pCf-ornU0b .VfPpkd-Bz112c-Jh9lGc::before,.jR8x9d .zF2sRd .VfPpkd-Cv7pCf-ornU0b .VfPpkd-Bz112c-Jh9lGc::after{background-color:rgb(232,234,237);background-color:var(--mdc-ripple-color,rgb(232,234,237))}.jR8x9d .zF2sRd .VfPpkd-Cv7pCf-ornU0b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.jR8x9d .zF2sRd .VfPpkd-Cv7pCf-ornU0b:not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(248,249,250)}.jR8x9d .zF2sRd .VfPpkd-Cv7pCf-ornU0b:not(:disabled):active{color:rgb(248,249,250)}.jR8x9d .zF2sRd.VfPpkd-Zc28rc-OWXEXe-xl07Ob-FNFY6c .VfPpkd-Cv7pCf-ornU0b{color:rgb(248,249,250);background-color:rgba(232,234,237,.12)}.jR8x9d .zF2sRd .VfPpkd-Cv7pCf-ornU0b:hover,.jR8x9d .zF2sRd .VfPpkd-oEZKA:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-Cv7pCf-ornU0b{color:rgb(248,249,250)}.jR8x9d .zF2sRd .VfPpkd-Cv7pCf-ornU0b:hover:disabled,.jR8x9d .zF2sRd .VfPpkd-oEZKA:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-Cv7pCf-ornU0b:disabled{color:rgba(232,234,237,.38)}.jR8x9d .cNUpL .VfPpkd-Cv7pCf-ornU0b{color:rgb(154,160,166)}.jR8x9d .cNUpL .VfPpkd-Cv7pCf-ornU0b:disabled{color:rgba(232,234,237,.38)}.jR8x9d .cNUpL .VfPpkd-Cv7pCf-ornU0b .VfPpkd-Bz112c-Jh9lGc::before,.jR8x9d .cNUpL .VfPpkd-Cv7pCf-ornU0b .VfPpkd-Bz112c-Jh9lGc::after{background-color:rgb(232,234,237);background-color:var(--mdc-ripple-color,rgb(232,234,237))}.jR8x9d .cNUpL .VfPpkd-Cv7pCf-ornU0b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.jR8x9d .cNUpL .VfPpkd-Cv7pCf-ornU0b:not(.VfPpkd-ksKsZd-mWPk3d):focus{color:rgb(248,249,250)}.jR8x9d .cNUpL .VfPpkd-Cv7pCf-ornU0b:not(:disabled):active{color:rgb(248,249,250)}.jR8x9d .cNUpL.VfPpkd-Zc28rc-OWXEXe-xl07Ob-FNFY6c .VfPpkd-Cv7pCf-ornU0b{color:rgb(248,249,250);background-color:rgba(232,234,237,.12)}.jR8x9d .cNUpL .VfPpkd-Cv7pCf-ornU0b:hover,.jR8x9d .cNUpL .VfPpkd-oEZKA:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-Cv7pCf-ornU0b{color:rgb(248,249,250)}.jR8x9d .cNUpL .VfPpkd-Cv7pCf-ornU0b:hover:disabled,.jR8x9d .cNUpL .VfPpkd-oEZKA:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-Cv7pCf-ornU0b:disabled{color:rgba(232,234,237,.38)}.jR8x9d .UDxLd .VfPpkd-k2Wrsb{color:#e8eaed}.jR8x9d .UDxLd .VfPpkd-cnG4Wd{color:#9aa0a6}.jR8x9d .UDxLd .VfPpkd-zMU9ub{color:rgb(154,160,166)}.jR8x9d .UDxLd .VfPpkd-zMU9ub .VfPpkd-Bz112c-Jh9lGc::before,.jR8x9d .UDxLd .VfPpkd-zMU9ub .VfPpkd-Bz112c-Jh9lGc::after{background-color:rgb(154,160,166);background-color:var(--mdc-ripple-color,rgb(154,160,166))}.jR8x9d .UDxLd .VfPpkd-zMU9ub:hover .VfPpkd-Bz112c-Jh9lGc::before,.jR8x9d .UDxLd .VfPpkd-zMU9ub.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Bz112c-Jh9lGc::before{opacity:.08;opacity:var(--mdc-ripple-hover-opacity,.08)}.jR8x9d .UDxLd .VfPpkd-zMU9ub.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Bz112c-Jh9lGc::before,.jR8x9d .UDxLd .VfPpkd-zMU9ub:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Bz112c-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.24;opacity:var(--mdc-ripple-focus-opacity,.24)}.jR8x9d .UDxLd .VfPpkd-zMU9ub:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Bz112c-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .UDxLd .VfPpkd-zMU9ub:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Bz112c-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.24;opacity:var(--mdc-ripple-press-opacity,.24)}.jR8x9d .UDxLd .VfPpkd-zMU9ub.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.24)}.jR8x9d .UDxLd .VfPpkd-IE5DDf,.jR8x9d .UDxLd .VfPpkd-P5QLlc-GGAcbc{background-color:rgba(0,0,0,.87)}.jR8x9d .UDxLd .VfPpkd-P5QLlc{background-color:rgb(32,33,36)}.jR8x9d .UDxLd .VfPpkd-P5QLlc{border-width:0;box-shadow:0 1px 3px 0 rgba(0,0,0,.3),0 4px 8px 3px rgba(0,0,0,.15)}.jR8x9d .UDxLd .VfPpkd-P5QLlc .VfPpkd-BFbNVe-bF1uUb{opacity:.11}.jR8x9d .ZD5Qo{color:rgb(138,180,248)}.jR8x9d .NNFoTc{background-color:rgb(32,33,36);height:56px;width:56px;padding-top:2px;padding-top:max(0px,2px);padding-right:2px;padding-right:max(0px,2px);padding-bottom:2px;padding-bottom:max(0px,2px);padding-left:2px;padding-left:max(0px,2px)}.jR8x9d .NNFoTc:not(:disabled){box-shadow:0 1px 3px 0 rgba(0,0,0,.3),0 4px 8px 3px rgba(0,0,0,.15)}.jR8x9d .NNFoTc:not(:disabled) .VfPpkd-BFbNVe-bF1uUb{opacity:.11}.jR8x9d .NNFoTc:not(:disabled) .VfPpkd-BFbNVe-bF1uUb{background-color:rgb(232,234,237)}.jR8x9d .NNFoTc:not(:disabled):hover{box-shadow:0 2px 3px 0 rgba(0,0,0,.3),0 6px 10px 4px rgba(0,0,0,.15)}.jR8x9d .NNFoTc:not(:disabled):hover .VfPpkd-BFbNVe-bF1uUb{opacity:.12}.jR8x9d .NNFoTc:not(:disabled):hover .VfPpkd-BFbNVe-bF1uUb{background-color:rgb(232,234,237)}.jR8x9d .NNFoTc:not(:disabled):focus{box-shadow:0 1px 3px 0 rgba(0,0,0,.3),0 4px 8px 3px rgba(0,0,0,.15)}.jR8x9d .NNFoTc:not(:disabled):focus .VfPpkd-BFbNVe-bF1uUb{opacity:.11}.jR8x9d .NNFoTc:not(:disabled):focus .VfPpkd-BFbNVe-bF1uUb{background-color:rgb(232,234,237)}.jR8x9d .NNFoTc:not(:disabled):active{box-shadow:0 4px 4px 0 rgba(0,0,0,.3),0 8px 12px 6px rgba(0,0,0,.15)}.jR8x9d .NNFoTc:not(:disabled):active .VfPpkd-BFbNVe-bF1uUb{opacity:.14}.jR8x9d .NNFoTc:not(:disabled):active .VfPpkd-BFbNVe-bF1uUb{background-color:rgb(232,234,237)}.jR8x9d .NNFoTc:disabled{box-shadow:0 1px 3px 0 rgba(0,0,0,.3),0 4px 8px 3px rgba(0,0,0,.15)}.jR8x9d .NNFoTc:disabled .VfPpkd-BFbNVe-bF1uUb{opacity:.11}.jR8x9d .NNFoTc:disabled .VfPpkd-BFbNVe-bF1uUb{background-color:rgb(232,234,237)}.jR8x9d .NNFoTc .VfPpkd-Q0XOV{width:36px;height:36px;font-size:36px}.jR8x9d .NNFoTc:not(:disabled) .VfPpkd-Q0XOV{color:rgb(232,234,237)}.jR8x9d .NNFoTc:not(:disabled):hover .VfPpkd-Q0XOV{color:rgb(174,203,250)}.jR8x9d .NNFoTc:not(:disabled):focus .VfPpkd-Q0XOV{color:rgb(174,203,250)}.jR8x9d .NNFoTc .VfPpkd-wbSZ0b::before,.jR8x9d .NNFoTc .VfPpkd-wbSZ0b::after{background-color:rgb(138,180,248)}.jR8x9d .NNFoTc:hover .VfPpkd-wbSZ0b::before,.jR8x9d .NNFoTc.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-wbSZ0b::before{opacity:.04}.jR8x9d .NNFoTc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-wbSZ0b::before,.jR8x9d .NNFoTc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-wbSZ0b::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12}.jR8x9d .NNFoTc:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-wbSZ0b::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .NNFoTc:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-wbSZ0b::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1}.jR8x9d .NNFoTc.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-fab-pressed-state-layer-opacity,0.1)}.jR8x9d .NNFoTc:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.jR8x9d .NNFoTc:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{border-color:rgb(102,157,246)}.jR8x9d .NNFoTc:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.jR8x9d .NNFoTc:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{border-style:solid;border-width:2px;padding-top:2px;padding-top:max(-2px,2px);padding-right:2px;padding-right:max(-2px,2px);padding-bottom:2px;padding-bottom:max(-2px,2px);padding-left:2px;padding-left:max(-2px,2px)}.jR8x9d .NNFoTc:not(.VfPpkd-BIzmGd-OWXEXe-X9G3K){border-radius:28px 28px 28px 28px}.jR8x9d .NNFoTc:not(.VfPpkd-BIzmGd-OWXEXe-X9G3K) .VfPpkd-wbSZ0b{border-radius:28px 28px 28px 28px}.jR8x9d .gl6QPb{background-color:rgb(32,33,36);height:48px;padding-top:max(0px,2px);padding-right:2px;padding-right:max(0px,2px);padding-bottom:max(0px,2px);padding-left:2px;padding-left:max(0px,2px);border-radius:24px 24px 24px 24px;font-family:Google Sans,Roboto,Arial,sans-serif;font-size:.875rem;font-weight:500;letter-spacing:.0178571429em;padding-top:2px;padding-right:24px;padding-bottom:2px;padding-left:24px}.jR8x9d .gl6QPb:not(:disabled){box-shadow:0 1px 3px 0 rgba(0,0,0,.3),0 4px 8px 3px rgba(0,0,0,.15)}.jR8x9d .gl6QPb:not(:disabled) .VfPpkd-BFbNVe-bF1uUb{opacity:.11}.jR8x9d .gl6QPb:not(:disabled) .VfPpkd-BFbNVe-bF1uUb{background-color:rgb(232,234,237)}.jR8x9d .gl6QPb:not(:disabled):hover{box-shadow:0 2px 3px 0 rgba(0,0,0,.3),0 6px 10px 4px rgba(0,0,0,.15)}.jR8x9d .gl6QPb:not(:disabled):hover .VfPpkd-BFbNVe-bF1uUb{opacity:.12}.jR8x9d .gl6QPb:not(:disabled):hover .VfPpkd-BFbNVe-bF1uUb{background-color:rgb(232,234,237)}.jR8x9d .gl6QPb:not(:disabled):focus{box-shadow:0 1px 3px 0 rgba(0,0,0,.3),0 4px 8px 3px rgba(0,0,0,.15)}.jR8x9d .gl6QPb:not(:disabled):focus .VfPpkd-BFbNVe-bF1uUb{opacity:.11}.jR8x9d .gl6QPb:not(:disabled):focus .VfPpkd-BFbNVe-bF1uUb{background-color:rgb(232,234,237)}.jR8x9d .gl6QPb:not(:disabled):active{box-shadow:0 4px 4px 0 rgba(0,0,0,.3),0 8px 12px 6px rgba(0,0,0,.15)}.jR8x9d .gl6QPb:not(:disabled):active .VfPpkd-BFbNVe-bF1uUb{opacity:.14}.jR8x9d .gl6QPb:not(:disabled):active .VfPpkd-BFbNVe-bF1uUb{background-color:rgb(232,234,237)}.jR8x9d .gl6QPb:disabled{box-shadow:0 1px 3px 0 rgba(0,0,0,.3),0 4px 8px 3px rgba(0,0,0,.15)}.jR8x9d .gl6QPb:disabled .VfPpkd-BFbNVe-bF1uUb{opacity:.11}.jR8x9d .gl6QPb:disabled .VfPpkd-BFbNVe-bF1uUb{background-color:rgb(232,234,237)}.jR8x9d .gl6QPb .VfPpkd-Q0XOV{width:36px;height:36px;font-size:36px}.jR8x9d .gl6QPb:not(:disabled) .VfPpkd-Q0XOV{color:rgb(232,234,237)}.jR8x9d .gl6QPb:not(:disabled):hover .VfPpkd-Q0XOV{color:rgb(174,203,250)}.jR8x9d .gl6QPb:not(:disabled):focus .VfPpkd-Q0XOV{color:rgb(174,203,250)}.jR8x9d .gl6QPb .VfPpkd-wbSZ0b::before,.jR8x9d .gl6QPb .VfPpkd-wbSZ0b::after{background-color:rgb(138,180,248)}.jR8x9d .gl6QPb:hover .VfPpkd-wbSZ0b::before,.jR8x9d .gl6QPb.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-wbSZ0b::before{opacity:.04}.jR8x9d .gl6QPb.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-wbSZ0b::before,.jR8x9d .gl6QPb:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-wbSZ0b::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12}.jR8x9d .gl6QPb:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-wbSZ0b::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .gl6QPb:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-wbSZ0b::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1}.jR8x9d .gl6QPb.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-extended-fab-pressed-state-layer-opacity,0.1)}.jR8x9d .gl6QPb:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.jR8x9d .gl6QPb:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{border-color:rgb(102,157,246)}.jR8x9d .gl6QPb:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.jR8x9d .gl6QPb:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{padding-top:max(-2px,2px);padding-right:2px;padding-right:max(-2px,2px);padding-bottom:max(-2px,2px);padding-left:2px;padding-left:max(-2px,2px)}.jR8x9d .gl6QPb .VfPpkd-wbSZ0b{border-radius:24px 24px 24px 24px}.jR8x9d .gl6QPb:not(:disabled) .VfPpkd-nBWOSb{color:rgb(232,234,237)}.jR8x9d .gl6QPb:not(:disabled):hover .VfPpkd-nBWOSb{color:rgb(174,203,250)}.jR8x9d .gl6QPb:not(:disabled):focus .VfPpkd-nBWOSb{color:rgb(174,203,250)}.jR8x9d .gl6QPb:not(:disabled):active .VfPpkd-nBWOSb{color:rgb(174,203,250)}.jR8x9d .gl6QPb .VfPpkd-Q0XOV{margin-left:-12px;margin-right:12px}[dir=rtl] .jR8x9d .gl6QPb .VfPpkd-Q0XOV,.jR8x9d .gl6QPb .VfPpkd-Q0XOV[dir=rtl]{margin-left:12px;margin-right:-12px}.jR8x9d .gl6QPb .VfPpkd-nBWOSb+.VfPpkd-Q0XOV{margin-left:12px;margin-right:-12px}[dir=rtl] .jR8x9d .gl6QPb .VfPpkd-nBWOSb+.VfPpkd-Q0XOV,.jR8x9d .gl6QPb .VfPpkd-nBWOSb+.VfPpkd-Q0XOV[dir=rtl]{margin-left:-12px;margin-right:12px}.jR8x9d .gl6QPb:not(:disabled).VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe,.jR8x9d .gl6QPb:not(:disabled):not(.VfPpkd-ksKsZd-mWPk3d):focus{border-style:solid;border-width:2px;padding-top:2px;padding-right:22px;padding-bottom:2px;padding-left:22px}.jR8x9d .Aykzec{background-color:rgb(138,180,248);height:48px;border-radius:24px 24px 24px 24px;font-family:Google Sans,Roboto,Arial,sans-serif;font-size:.875rem;font-weight:500;letter-spacing:.0178571429em}.jR8x9d .Aykzec:not(:disabled){box-shadow:0 1px 3px 0 rgba(0,0,0,.3),0 4px 8px 3px rgba(0,0,0,.15)}.jR8x9d .Aykzec:not(:disabled) .VfPpkd-BFbNVe-bF1uUb{opacity:.11}.jR8x9d .Aykzec:not(:disabled) .VfPpkd-BFbNVe-bF1uUb{background-color:rgb(232,234,237)}.jR8x9d .Aykzec:not(:disabled):hover{box-shadow:0 2px 3px 0 rgba(0,0,0,.3),0 6px 10px 4px rgba(0,0,0,.15)}.jR8x9d .Aykzec:not(:disabled):hover .VfPpkd-BFbNVe-bF1uUb{opacity:.12}.jR8x9d .Aykzec:not(:disabled):hover .VfPpkd-BFbNVe-bF1uUb{background-color:rgb(232,234,237)}.jR8x9d .Aykzec:not(:disabled):focus{box-shadow:0 1px 3px 0 rgba(0,0,0,.3),0 4px 8px 3px rgba(0,0,0,.15)}.jR8x9d .Aykzec:not(:disabled):focus .VfPpkd-BFbNVe-bF1uUb{opacity:.11}.jR8x9d .Aykzec:not(:disabled):focus .VfPpkd-BFbNVe-bF1uUb{background-color:rgb(232,234,237)}.jR8x9d .Aykzec:not(:disabled):active{box-shadow:0 4px 4px 0 rgba(0,0,0,.3),0 8px 12px 6px rgba(0,0,0,.15)}.jR8x9d .Aykzec:not(:disabled):active .VfPpkd-BFbNVe-bF1uUb{opacity:.14}.jR8x9d .Aykzec:not(:disabled):active .VfPpkd-BFbNVe-bF1uUb{background-color:rgb(232,234,237)}.jR8x9d .Aykzec:disabled{box-shadow:0 1px 3px 0 rgba(0,0,0,.3),0 4px 8px 3px rgba(0,0,0,.15)}.jR8x9d .Aykzec:disabled .VfPpkd-BFbNVe-bF1uUb{opacity:.11}.jR8x9d .Aykzec:disabled .VfPpkd-BFbNVe-bF1uUb{background-color:rgb(232,234,237)}.jR8x9d .Aykzec .VfPpkd-Q0XOV{width:24px;height:24px;font-size:24px}.jR8x9d .Aykzec:not(:disabled) .VfPpkd-Q0XOV{color:rgb(32,33,36)}.jR8x9d .Aykzec .VfPpkd-wbSZ0b::before,.jR8x9d .Aykzec .VfPpkd-wbSZ0b::after{background-color:rgb(255,255,255)}.jR8x9d .Aykzec:hover .VfPpkd-wbSZ0b::before,.jR8x9d .Aykzec.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-wbSZ0b::before{opacity:.16}.jR8x9d .Aykzec.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-wbSZ0b::before,.jR8x9d .Aykzec:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-wbSZ0b::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.24}.jR8x9d .Aykzec:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-wbSZ0b::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .Aykzec:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-wbSZ0b::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.2}.jR8x9d .Aykzec.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-extended-fab-pressed-state-layer-opacity,0.2)}.jR8x9d .Aykzec .VfPpkd-wbSZ0b{border-radius:24px 24px 24px 24px}.jR8x9d .Aykzec:not(:disabled) .VfPpkd-nBWOSb{color:rgb(32,33,36)}.jR8x9d .W7mYUe{background-color:rgb(32,33,36);height:48px;border-radius:24px 24px 24px 24px;font-family:Google Sans,Roboto,Arial,sans-serif;font-size:.875rem;font-weight:500;letter-spacing:.0178571429em}.jR8x9d .W7mYUe:not(:disabled){box-shadow:0 1px 3px 0 rgba(0,0,0,.3),0 4px 8px 3px rgba(0,0,0,.15)}.jR8x9d .W7mYUe:not(:disabled) .VfPpkd-BFbNVe-bF1uUb{opacity:.11}.jR8x9d .W7mYUe:not(:disabled) .VfPpkd-BFbNVe-bF1uUb{background-color:rgb(232,234,237)}.jR8x9d .W7mYUe:not(:disabled):hover{box-shadow:0 2px 3px 0 rgba(0,0,0,.3),0 6px 10px 4px rgba(0,0,0,.15)}.jR8x9d .W7mYUe:not(:disabled):hover .VfPpkd-BFbNVe-bF1uUb{opacity:.12}.jR8x9d .W7mYUe:not(:disabled):hover .VfPpkd-BFbNVe-bF1uUb{background-color:rgb(232,234,237)}.jR8x9d .W7mYUe:not(:disabled):focus{box-shadow:0 1px 3px 0 rgba(0,0,0,.3),0 4px 8px 3px rgba(0,0,0,.15)}.jR8x9d .W7mYUe:not(:disabled):focus .VfPpkd-BFbNVe-bF1uUb{opacity:.11}.jR8x9d .W7mYUe:not(:disabled):focus .VfPpkd-BFbNVe-bF1uUb{background-color:rgb(232,234,237)}.jR8x9d .W7mYUe:not(:disabled):active{box-shadow:0 4px 4px 0 rgba(0,0,0,.3),0 8px 12px 6px rgba(0,0,0,.15)}.jR8x9d .W7mYUe:not(:disabled):active .VfPpkd-BFbNVe-bF1uUb{opacity:.14}.jR8x9d .W7mYUe:not(:disabled):active .VfPpkd-BFbNVe-bF1uUb{background-color:rgb(232,234,237)}.jR8x9d .W7mYUe:disabled{box-shadow:0 1px 3px 0 rgba(0,0,0,.3),0 4px 8px 3px rgba(0,0,0,.15)}.jR8x9d .W7mYUe:disabled .VfPpkd-BFbNVe-bF1uUb{opacity:.11}.jR8x9d .W7mYUe:disabled .VfPpkd-BFbNVe-bF1uUb{background-color:rgb(232,234,237)}.jR8x9d .W7mYUe .VfPpkd-Q0XOV{width:24px;height:24px;font-size:24px}.jR8x9d .W7mYUe:not(:disabled) .VfPpkd-Q0XOV{color:rgb(138,180,248)}.jR8x9d .W7mYUe:not(:disabled):hover .VfPpkd-Q0XOV{color:rgb(174,203,250)}.jR8x9d .W7mYUe:not(:disabled):focus .VfPpkd-Q0XOV{color:rgb(174,203,250)}.jR8x9d .W7mYUe:not(:disabled):active .VfPpkd-Q0XOV{color:rgb(174,203,250)}.jR8x9d .W7mYUe .VfPpkd-wbSZ0b::before,.jR8x9d .W7mYUe .VfPpkd-wbSZ0b::after{background-color:rgb(138,180,248)}.jR8x9d .W7mYUe:hover .VfPpkd-wbSZ0b::before,.jR8x9d .W7mYUe.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-wbSZ0b::before{opacity:.04}.jR8x9d .W7mYUe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-wbSZ0b::before,.jR8x9d .W7mYUe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-wbSZ0b::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12}.jR8x9d .W7mYUe:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-wbSZ0b::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .W7mYUe:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-wbSZ0b::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1}.jR8x9d .W7mYUe.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-extended-fab-pressed-state-layer-opacity,0.1)}.jR8x9d .W7mYUe .VfPpkd-wbSZ0b{border-radius:24px 24px 24px 24px}.jR8x9d .W7mYUe:not(:disabled) .VfPpkd-nBWOSb{color:rgb(138,180,248)}.jR8x9d .W7mYUe:not(:disabled):hover .VfPpkd-nBWOSb{color:rgb(174,203,250)}.jR8x9d .W7mYUe:not(:disabled):focus .VfPpkd-nBWOSb{color:rgb(174,203,250)}.jR8x9d .W7mYUe:not(:disabled):active .VfPpkd-nBWOSb{color:rgb(174,203,250)}.jR8x9d .OoEosd{background-color:rgb(32,33,36);height:56px;width:56px}.jR8x9d .OoEosd:not(:disabled){box-shadow:0 1px 3px 0 rgba(0,0,0,.3),0 4px 8px 3px rgba(0,0,0,.15)}.jR8x9d .OoEosd:not(:disabled) .VfPpkd-BFbNVe-bF1uUb{opacity:.11}.jR8x9d .OoEosd:not(:disabled) .VfPpkd-BFbNVe-bF1uUb{background-color:rgb(232,234,237)}.jR8x9d .OoEosd:not(:disabled):hover{box-shadow:0 2px 3px 0 rgba(0,0,0,.3),0 6px 10px 4px rgba(0,0,0,.15)}.jR8x9d .OoEosd:not(:disabled):hover .VfPpkd-BFbNVe-bF1uUb{opacity:.12}.jR8x9d .OoEosd:not(:disabled):hover .VfPpkd-BFbNVe-bF1uUb{background-color:rgb(232,234,237)}.jR8x9d .OoEosd:not(:disabled):focus{box-shadow:0 1px 3px 0 rgba(0,0,0,.3),0 4px 8px 3px rgba(0,0,0,.15)}.jR8x9d .OoEosd:not(:disabled):focus .VfPpkd-BFbNVe-bF1uUb{opacity:.11}.jR8x9d .OoEosd:not(:disabled):focus .VfPpkd-BFbNVe-bF1uUb{background-color:rgb(232,234,237)}.jR8x9d .OoEosd:not(:disabled):active{box-shadow:0 4px 4px 0 rgba(0,0,0,.3),0 8px 12px 6px rgba(0,0,0,.15)}.jR8x9d .OoEosd:not(:disabled):active .VfPpkd-BFbNVe-bF1uUb{opacity:.14}.jR8x9d .OoEosd:not(:disabled):active .VfPpkd-BFbNVe-bF1uUb{background-color:rgb(232,234,237)}.jR8x9d .OoEosd:disabled{box-shadow:0 1px 3px 0 rgba(0,0,0,.3),0 4px 8px 3px rgba(0,0,0,.15)}.jR8x9d .OoEosd:disabled .VfPpkd-BFbNVe-bF1uUb{opacity:.11}.jR8x9d .OoEosd:disabled .VfPpkd-BFbNVe-bF1uUb{background-color:rgb(232,234,237)}.jR8x9d .OoEosd .VfPpkd-Q0XOV{width:24px;height:24px;font-size:24px}.jR8x9d .OoEosd:not(:disabled) .VfPpkd-Q0XOV{color:rgb(138,180,248)}.jR8x9d .OoEosd:not(:disabled):hover .VfPpkd-Q0XOV{color:rgb(174,203,250)}.jR8x9d .OoEosd:not(:disabled):focus .VfPpkd-Q0XOV{color:rgb(174,203,250)}.jR8x9d .OoEosd:not(:disabled):active .VfPpkd-Q0XOV{color:rgb(174,203,250)}.jR8x9d .OoEosd .VfPpkd-wbSZ0b::before,.jR8x9d .OoEosd .VfPpkd-wbSZ0b::after{background-color:rgb(138,180,248)}.jR8x9d .OoEosd:hover .VfPpkd-wbSZ0b::before,.jR8x9d .OoEosd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-wbSZ0b::before{opacity:.04}.jR8x9d .OoEosd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-wbSZ0b::before,.jR8x9d .OoEosd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-wbSZ0b::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12}.jR8x9d .OoEosd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-wbSZ0b::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .OoEosd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-wbSZ0b::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1}.jR8x9d .OoEosd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-fab-pressed-state-layer-opacity,0.1)}.jR8x9d .OoEosd:not(.VfPpkd-BIzmGd-OWXEXe-X9G3K){border-radius:28px 28px 28px 28px}.jR8x9d .OoEosd:not(.VfPpkd-BIzmGd-OWXEXe-X9G3K) .VfPpkd-wbSZ0b{border-radius:28px 28px 28px 28px}.jR8x9d .vd3sk:not(:disabled){box-shadow:0 1px 2px 0 rgba(0,0,0,.3),0 1px 3px 1px rgba(0,0,0,.15)}.jR8x9d .vd3sk:not(:disabled) .VfPpkd-BFbNVe-bF1uUb{opacity:.05}.jR8x9d .vd3sk:not(:disabled) .VfPpkd-BFbNVe-bF1uUb{background-color:rgb(232,234,237)}.jR8x9d .vd3sk:not(:disabled):hover{box-shadow:0 1px 2px 0 rgba(0,0,0,.3),0 2px 6px 2px rgba(0,0,0,.15)}.jR8x9d .vd3sk:not(:disabled):hover .VfPpkd-BFbNVe-bF1uUb{opacity:.08}.jR8x9d .vd3sk:not(:disabled):hover .VfPpkd-BFbNVe-bF1uUb{background-color:rgb(232,234,237)}.jR8x9d .vd3sk:not(:disabled):focus{box-shadow:0 1px 2px 0 rgba(0,0,0,.3),0 2px 6px 2px rgba(0,0,0,.15)}.jR8x9d .vd3sk:not(:disabled):focus .VfPpkd-BFbNVe-bF1uUb{opacity:.08}.jR8x9d .vd3sk:not(:disabled):focus .VfPpkd-BFbNVe-bF1uUb{background-color:rgb(232,234,237)}.jR8x9d .vd3sk:not(:disabled):active{box-shadow:0 1px 3px 0 rgba(0,0,0,.3),0 4px 8px 3px rgba(0,0,0,.15)}.jR8x9d .vd3sk:not(:disabled):active .VfPpkd-BFbNVe-bF1uUb{opacity:.11}.jR8x9d .vd3sk:not(:disabled):active .VfPpkd-BFbNVe-bF1uUb{background-color:rgb(232,234,237)}.jR8x9d .vd3sk:disabled{box-shadow:0 1px 2px 0 rgba(0,0,0,.3),0 1px 3px 1px rgba(0,0,0,.15)}.jR8x9d .vd3sk:disabled .VfPpkd-BFbNVe-bF1uUb{opacity:.05}.jR8x9d .vd3sk:disabled .VfPpkd-BFbNVe-bF1uUb{background-color:rgb(232,234,237)}.jR8x9d .N7pe4e:not(:disabled){box-shadow:0 1px 2px 0 rgba(0,0,0,.3),0 1px 3px 1px rgba(0,0,0,.15)}.jR8x9d .N7pe4e:not(:disabled) .VfPpkd-BFbNVe-bF1uUb{opacity:.05}.jR8x9d .N7pe4e:not(:disabled) .VfPpkd-BFbNVe-bF1uUb{background-color:rgb(232,234,237)}.jR8x9d .N7pe4e:not(:disabled):hover{box-shadow:0 1px 2px 0 rgba(0,0,0,.3),0 2px 6px 2px rgba(0,0,0,.15)}.jR8x9d .N7pe4e:not(:disabled):hover .VfPpkd-BFbNVe-bF1uUb{opacity:.08}.jR8x9d .N7pe4e:not(:disabled):hover .VfPpkd-BFbNVe-bF1uUb{background-color:rgb(232,234,237)}.jR8x9d .N7pe4e:not(:disabled):focus{box-shadow:0 1px 2px 0 rgba(0,0,0,.3),0 2px 6px 2px rgba(0,0,0,.15)}.jR8x9d .N7pe4e:not(:disabled):focus .VfPpkd-BFbNVe-bF1uUb{opacity:.08}.jR8x9d .N7pe4e:not(:disabled):focus .VfPpkd-BFbNVe-bF1uUb{background-color:rgb(232,234,237)}.jR8x9d .N7pe4e:not(:disabled):active{box-shadow:0 1px 3px 0 rgba(0,0,0,.3),0 4px 8px 3px rgba(0,0,0,.15)}.jR8x9d .N7pe4e:not(:disabled):active .VfPpkd-BFbNVe-bF1uUb{opacity:.11}.jR8x9d .N7pe4e:not(:disabled):active .VfPpkd-BFbNVe-bF1uUb{background-color:rgb(232,234,237)}.jR8x9d .N7pe4e:disabled{box-shadow:0 1px 2px 0 rgba(0,0,0,.3),0 1px 3px 1px rgba(0,0,0,.15)}.jR8x9d .N7pe4e:disabled .VfPpkd-BFbNVe-bF1uUb{opacity:.05}.jR8x9d .N7pe4e:disabled .VfPpkd-BFbNVe-bF1uUb{background-color:rgb(232,234,237)}.jR8x9d .JJMOVe:not(:disabled){box-shadow:0 1px 2px 0 rgba(0,0,0,.3),0 1px 3px 1px rgba(0,0,0,.15)}.jR8x9d .JJMOVe:not(:disabled) .VfPpkd-BFbNVe-bF1uUb{opacity:.05}.jR8x9d .JJMOVe:not(:disabled) .VfPpkd-BFbNVe-bF1uUb{background-color:rgb(232,234,237)}.jR8x9d .JJMOVe:not(:disabled):hover{box-shadow:0 1px 2px 0 rgba(0,0,0,.3),0 2px 6px 2px rgba(0,0,0,.15)}.jR8x9d .JJMOVe:not(:disabled):hover .VfPpkd-BFbNVe-bF1uUb{opacity:.08}.jR8x9d .JJMOVe:not(:disabled):hover .VfPpkd-BFbNVe-bF1uUb{background-color:rgb(232,234,237)}.jR8x9d .JJMOVe:not(:disabled):focus{box-shadow:0 1px 2px 0 rgba(0,0,0,.3),0 2px 6px 2px rgba(0,0,0,.15)}.jR8x9d .JJMOVe:not(:disabled):focus .VfPpkd-BFbNVe-bF1uUb{opacity:.08}.jR8x9d .JJMOVe:not(:disabled):focus .VfPpkd-BFbNVe-bF1uUb{background-color:rgb(232,234,237)}.jR8x9d .JJMOVe:not(:disabled):active{box-shadow:0 1px 3px 0 rgba(0,0,0,.3),0 4px 8px 3px rgba(0,0,0,.15)}.jR8x9d .JJMOVe:not(:disabled):active .VfPpkd-BFbNVe-bF1uUb{opacity:.11}.jR8x9d .JJMOVe:not(:disabled):active .VfPpkd-BFbNVe-bF1uUb{background-color:rgb(232,234,237)}.jR8x9d .JJMOVe:disabled{box-shadow:0 1px 2px 0 rgba(0,0,0,.3),0 1px 3px 1px rgba(0,0,0,.15)}.jR8x9d .JJMOVe:disabled .VfPpkd-BFbNVe-bF1uUb{opacity:.05}.jR8x9d .JJMOVe:disabled .VfPpkd-BFbNVe-bF1uUb{background-color:rgb(232,234,237)}.jR8x9d .E9mvxc{height:40px;width:40px}.jR8x9d .ZCuY4{font-family:Roboto,Arial,sans-serif;line-height:1.25rem;font-size:.875rem;letter-spacing:.0142857143em;font-weight:400;color:rgb(232,234,237)}.jR8x9d .ZCuY4 gm-checkbox[disabled]~.VfPpkd-V67aGc,.jR8x9d .ZCuY4 gm-radio[disabled]~.VfPpkd-V67aGc,.jR8x9d .ZCuY4 .VfPpkd-MPu53c-OWXEXe-OWB6Me~.VfPpkd-V67aGc,.jR8x9d .ZCuY4 .VfPpkd-GCYh9b-OWXEXe-OWB6Me~.VfPpkd-V67aGc{color:rgba(232,234,237,.38)}.jR8x9d .E2obDf .VfPpkd-qNpTzb-P4pF8c-SmKAyb{border-color:rgb(102,157,246)}.jR8x9d .E2obDf .VfPpkd-qNpTzb-ajuXxc-RxYbNe{background-color:rgba(138,180,248,.24)}}@media screen and (prefers-color-scheme:dark) and (forced-colors:active){.jR8x9d .E2obDf .VfPpkd-qNpTzb-ajuXxc-RxYbNe{background-color:ButtonBorder}}@media screen and (prefers-color-scheme:dark) and (-ms-high-contrast:active),screen and (prefers-color-scheme:dark) and (-ms-high-contrast:none){.jR8x9d .E2obDf .VfPpkd-qNpTzb-ajuXxc-RxYbNe{background-color:transparent;background-image:url("data:image/svg+xml,%3Csvg version='1.1' xmlns='http://www.w3.org/2000/svg' xmlns:xlink='http://www.w3.org/1999/xlink' x='0px' y='0px' enable-background='new 0 0 5 2' xml:space='preserve' viewBox='0 0 5 2' preserveAspectRatio='none slice'%3E%3Ccircle cx='1' cy='1' r='1' fill='rgba(138, 180, 248, 0.24)'/%3E%3C/svg%3E")}}@media screen and (prefers-color-scheme:dark){.jR8x9d .E2obDf .VfPpkd-qNpTzb-ajuXxc-ZMv3u{background-color:rgba(138,180,248,.24)}.jR8x9d .bwNLcf{color:rgb(232,234,237);font-family:Roboto,Arial,sans-serif;line-height:1.5rem;font-size:1rem;letter-spacing:.00625em;font-weight:400}.jR8x9d .bwNLcf .VfPpkd-StrnGf-rymPhb-IhFlZd{color:rgb(154,160,166)}.jR8x9d .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.jR8x9d .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.jR8x9d .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS{color:rgb(232,234,237)}.jR8x9d .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c{opacity:.38}.jR8x9d .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd,.jR8x9d .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b,.jR8x9d .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-f7MjDc,.jR8x9d .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-f7MjDc{color:rgb(232,234,237)}.jR8x9d .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:0}.jR8x9d .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd{background-color:rgba(138,180,248,.24)}.jR8x9d .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before,.jR8x9d .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::after{background-color:rgb(138,180,248);background-color:var(--mdc-ripple-color,rgb(138,180,248))}.jR8x9d .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before,.jR8x9d .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.jR8x9d .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before,.jR8x9d .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.jR8x9d .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.jR8x9d .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}.jR8x9d .bwNLcf .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS{color:rgb(154,160,166)}.jR8x9d .bwNLcf .VfPpkd-StrnGf-rymPhb-clz4Ic{border-bottom-color:rgba(232,234,237,.12)}.jR8x9d .bwNLcf .VfPpkd-StrnGf-rymPhb-f7MjDc{color:rgb(232,234,237)}.jR8x9d .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-pZXsl::before,.jR8x9d .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-pZXsl::after{background-color:rgb(232,234,237);background-color:var(--mdc-ripple-color,rgb(232,234,237))}.jR8x9d .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before,.jR8x9d .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.jR8x9d .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before,.jR8x9d .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.jR8x9d .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.jR8x9d .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}}@media screen and (prefers-color-scheme:dark) and (-ms-high-contrast:active),screen and (prefers-color-scheme:dark) and (forced-colors:active){.jR8x9d .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.jR8x9d .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.jR8x9d .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS{color:GrayText}.jR8x9d .bwNLcf .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c{opacity:1}}@media screen and (prefers-color-scheme:dark){.jR8x9d .bwNLcf .VfPpkd-rymPhb-Gtdoyb,.jR8x9d .bwNLcf .VfPpkd-rymPhb-fpDzbe-fmcmS{color:rgb(232,234,237)}.jR8x9d .bwNLcf .VfPpkd-rymPhb-L8ivfd-fmcmS,.jR8x9d .bwNLcf .VfPpkd-rymPhb-bC5pod-fmcmS,.jR8x9d .bwNLcf .VfPpkd-rymPhb-JMEf7e{color:rgb(154,160,166)}.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb,.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e,.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-Gtdoyb,.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-fpDzbe-fmcmS,.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-L8ivfd-fmcmS,.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-bC5pod-fmcmS,.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb,.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e,.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e{color:rgb(232,234,237)}.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-KkROqb,.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-Gtdoyb,.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-JMEf7e{opacity:.38}.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-Gtdoyb,.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-fpDzbe-fmcmS,.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-rymPhb-Gtdoyb,.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-rymPhb-fpDzbe-fmcmS,.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb,.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb{color:rgb(232,234,237)}.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::before{opacity:0}.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd{background-color:rgba(138,180,248,.24)}.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::before,.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::after{background-color:rgb(138,180,248);background-color:var(--mdc-ripple-color,rgb(138,180,248))}.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-rymPhb-pZXsl::before,.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-rymPhb-pZXsl::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-rymPhb-pZXsl::before,.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-rymPhb-pZXsl::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-rymPhb-pZXsl::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-rymPhb-pZXsl::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}.jR8x9d .bwNLcf .VfPpkd-rymPhb-L8ivfd-fmcmS{color:rgb(154,160,166)}.jR8x9d .bwNLcf .VfPpkd-rymPhb-clz4Ic{background-color:rgba(232,234,237,.12)}.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb,.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e{color:rgb(232,234,237)}.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::before,.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::after{background-color:rgb(232,234,237);background-color:var(--mdc-ripple-color,rgb(232,234,237))}.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b:hover .VfPpkd-rymPhb-pZXsl::before,.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-rymPhb-pZXsl::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-rymPhb-pZXsl::before,.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-rymPhb-pZXsl::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-rymPhb-pZXsl::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-rymPhb-pZXsl::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}}@media screen and (prefers-color-scheme:dark) and (forced-colors:active){.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-Gtdoyb,.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-fpDzbe-fmcmS,.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-L8ivfd-fmcmS,.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-bC5pod-fmcmS,.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb,.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e,.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e{color:GrayText}.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-KkROqb,.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-Gtdoyb,.jR8x9d .bwNLcf .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-JMEf7e{opacity:1}}@media screen and (prefers-color-scheme:dark){.jR8x9d .f8F5Dd{background-color:rgb(32,33,36);border-width:0;box-shadow:0 1px 2px 0 rgba(0,0,0,.3),0 2px 6px 2px rgba(0,0,0,.15)}.jR8x9d .f8F5Dd .VfPpkd-BFbNVe-bF1uUb{opacity:.08}.jR8x9d .P77izf{background-color:rgb(32,33,36);border-width:0;box-shadow:0 1px 2px 0 rgba(0,0,0,.3),0 2px 6px 2px rgba(0,0,0,.15)}.jR8x9d .P77izf .VfPpkd-StrnGf-rymPhb{font-family:Roboto,Arial,sans-serif;line-height:1.5rem;font-size:1rem;letter-spacing:.00625em;font-weight:400;color:rgb(232,234,237)}.jR8x9d .P77izf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-IhFlZd{color:rgb(154,160,166)}.jR8x9d .P77izf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.jR8x9d .P77izf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.jR8x9d .P77izf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS{color:rgb(232,234,237)}.jR8x9d .P77izf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c{opacity:.38}.jR8x9d .P77izf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd,.jR8x9d .P77izf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b,.jR8x9d .P77izf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-f7MjDc,.jR8x9d .P77izf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-f7MjDc{color:rgb(232,234,237)}.jR8x9d .P77izf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:0}.jR8x9d .P77izf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd{background-color:rgba(138,180,248,.24)}.jR8x9d .P77izf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before,.jR8x9d .P77izf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::after{background-color:rgb(138,180,248);background-color:var(--mdc-ripple-color,rgb(138,180,248))}.jR8x9d .P77izf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before,.jR8x9d .P77izf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.jR8x9d .P77izf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before,.jR8x9d .P77izf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.jR8x9d .P77izf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .P77izf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.jR8x9d .P77izf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}.jR8x9d .P77izf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS{color:rgb(154,160,166)}.jR8x9d .P77izf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic{border-bottom-color:rgba(232,234,237,.12)}.jR8x9d .P77izf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc{color:rgb(232,234,237)}.jR8x9d .P77izf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-pZXsl::before,.jR8x9d .P77izf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-pZXsl::after{background-color:rgb(232,234,237);background-color:var(--mdc-ripple-color,rgb(232,234,237))}.jR8x9d .P77izf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before,.jR8x9d .P77izf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.jR8x9d .P77izf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before,.jR8x9d .P77izf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.jR8x9d .P77izf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .P77izf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.jR8x9d .P77izf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}}@media screen and (prefers-color-scheme:dark) and (-ms-high-contrast:active),screen and (prefers-color-scheme:dark) and (forced-colors:active){.jR8x9d .P77izf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.jR8x9d .P77izf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.jR8x9d .P77izf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS{color:GrayText}.jR8x9d .P77izf .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c{opacity:1}}@media screen and (prefers-color-scheme:dark){.jR8x9d .P77izf .VfPpkd-BFbNVe-bF1uUb{opacity:.08}.jR8x9d .ZCYEwf{z-index:0}.jR8x9d .ZCYEwf .VfPpkd-eHTEvd::before,.jR8x9d .ZCYEwf .VfPpkd-eHTEvd::after{z-index:-1}.jR8x9d .ZCYEwf .VfPpkd-eHTEvd::before,.jR8x9d .ZCYEwf .VfPpkd-eHTEvd::after{background-color:rgb(138,180,248);background-color:var(--gm-radio-state-color,rgb(138,180,248))}.jR8x9d .ZCYEwf:hover .VfPpkd-eHTEvd::before,.jR8x9d .ZCYEwf.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-eHTEvd::before{opacity:.16;opacity:var(--mdc-ripple-hover-opacity,.16)}.jR8x9d .ZCYEwf.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-eHTEvd::before,.jR8x9d .ZCYEwf:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-eHTEvd::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.24;opacity:var(--mdc-ripple-focus-opacity,.24)}.jR8x9d .ZCYEwf:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-eHTEvd::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .ZCYEwf:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-eHTEvd::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.2;opacity:var(--mdc-ripple-press-opacity,.2)}.jR8x9d .ZCYEwf .VfPpkd-gBXA9-bMcfAe:enabled:not(:checked)~.VfPpkd-eHTEvd::before,.jR8x9d .ZCYEwf .VfPpkd-gBXA9-bMcfAe:enabled:not(:checked)~.VfPpkd-eHTEvd::after{background-color:rgb(232,234,237);background-color:var(--gm-radio-state-color,rgb(232,234,237))}.jR8x9d .ZCYEwf:hover .VfPpkd-gBXA9-bMcfAe:enabled:not(:checked)~.VfPpkd-eHTEvd::before,.jR8x9d .ZCYEwf.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-gBXA9-bMcfAe:enabled:not(:checked)~.VfPpkd-eHTEvd::before{opacity:.16;opacity:var(--mdc-ripple-hover-opacity,.16)}.jR8x9d .ZCYEwf.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-gBXA9-bMcfAe:enabled:not(:checked)~.VfPpkd-eHTEvd::before,.jR8x9d .ZCYEwf:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-gBXA9-bMcfAe:enabled:not(:checked)~.VfPpkd-eHTEvd::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.24;opacity:var(--mdc-ripple-focus-opacity,.24)}.jR8x9d .ZCYEwf:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-gBXA9-bMcfAe:enabled:not(:checked)~.VfPpkd-eHTEvd::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .ZCYEwf:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-gBXA9-bMcfAe:enabled:not(:checked)~.VfPpkd-eHTEvd::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.2;opacity:var(--mdc-ripple-press-opacity,.2)}.jR8x9d .ZCYEwf.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.2)}.jR8x9d .ZCYEwf .VfPpkd-gBXA9-bMcfAe:enabled:not(:checked)+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgb(154,160,166);border-color:var(--gm-radio-stroke-color--unchecked,rgb(154,160,166))}.jR8x9d .ZCYEwf .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgb(138,180,248);border-color:var(--gm-radio-stroke-color--checked,rgb(138,180,248))}.jR8x9d .ZCYEwf .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo{border-color:rgb(138,180,248);border-color:var(--gm-radio-ink-color,rgb(138,180,248))}.jR8x9d .ZCYEwf [aria-disabled=true] .VfPpkd-gBXA9-bMcfAe:not(:checked)+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo,.jR8x9d .ZCYEwf .VfPpkd-gBXA9-bMcfAe:disabled:not(:checked)+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgba(232,234,237,.38);border-color:var(--gm-radio-disabled-stroke-color--unchecked,rgba(232,234,237,.38))}.jR8x9d .ZCYEwf [aria-disabled=true] .VfPpkd-gBXA9-bMcfAe:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo,.jR8x9d .ZCYEwf .VfPpkd-gBXA9-bMcfAe:disabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgba(232,234,237,.38);border-color:var(--gm-radio-disabled-stroke-color--checked,rgba(232,234,237,.38))}.jR8x9d .ZCYEwf [aria-disabled=true] .VfPpkd-gBXA9-bMcfAe+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo,.jR8x9d .ZCYEwf .VfPpkd-gBXA9-bMcfAe:disabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo{border-color:rgba(232,234,237,.38);border-color:var(--gm-radio-disabled-ink-color,rgba(232,234,237,.38))}.jR8x9d .ZCYEwf .VfPpkd-RsCWK::before{background-color:rgb(138,180,248);background-color:var(--gm-radio-state-color,rgb(138,180,248))}.jR8x9d .ZCYEwf:hover .VfPpkd-gBXA9-bMcfAe:enabled:not(:checked)+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo,.jR8x9d .ZCYEwf.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-gBXA9-bMcfAe:enabled:not(:checked)+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo,.jR8x9d .ZCYEwf:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-gBXA9-bMcfAe:enabled:not(:checked)+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo,.jR8x9d .ZCYEwf:active .VfPpkd-gBXA9-bMcfAe:enabled:not(:checked)+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgb(232,234,237);border-color:var(--gm-radio-stroke-color--unchecked-stateful,rgb(232,234,237))}.jR8x9d .ZCYEwf:hover .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo,.jR8x9d .ZCYEwf.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo,.jR8x9d .ZCYEwf:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo,.jR8x9d .ZCYEwf:active .VfPpkd-gBXA9-bMcfAe:enabled:checked+.VfPpkd-RsCWK .VfPpkd-wVo5xe-LkdAo{border-color:rgb(174,203,250);border-color:var(--gm-radio-stroke-color--checked-stateful,rgb(174,203,250))}.jR8x9d .ZCYEwf:hover .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo,.jR8x9d .ZCYEwf.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo,.jR8x9d .ZCYEwf:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo,.jR8x9d .ZCYEwf:active .VfPpkd-gBXA9-bMcfAe:enabled+.VfPpkd-RsCWK .VfPpkd-Z5TpLc-LkdAo{border-color:rgb(174,203,250);border-color:var(--gm-radio-ink-color--stateful,rgb(174,203,250))}.jR8x9d .dmaMHc{background-color:rgb(32,33,36);border-width:0;box-shadow:0 1px 2px 0 rgba(0,0,0,.3),0 2px 6px 2px rgba(0,0,0,.15);font-family:Roboto,Arial,sans-serif;line-height:1.5rem;font-size:1rem;letter-spacing:.00625em;font-weight:400}.jR8x9d .dmaMHc .VfPpkd-StrnGf-rymPhb{font-family:Roboto,Arial,sans-serif;line-height:1.5rem;font-size:1rem;letter-spacing:.00625em;font-weight:400;color:rgb(232,234,237)}.jR8x9d .dmaMHc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-IhFlZd{color:rgb(154,160,166)}.jR8x9d .dmaMHc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.jR8x9d .dmaMHc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.jR8x9d .dmaMHc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS{color:rgb(232,234,237)}.jR8x9d .dmaMHc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c{opacity:.38}.jR8x9d .dmaMHc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd,.jR8x9d .dmaMHc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b,.jR8x9d .dmaMHc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-f7MjDc,.jR8x9d .dmaMHc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-StrnGf-rymPhb-f7MjDc{color:rgb(232,234,237)}.jR8x9d .dmaMHc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:0}.jR8x9d .dmaMHc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd{background-color:rgba(138,180,248,.24)}.jR8x9d .dmaMHc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before,.jR8x9d .dmaMHc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::after{background-color:rgb(138,180,248);background-color:var(--mdc-ripple-color,rgb(138,180,248))}.jR8x9d .dmaMHc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before,.jR8x9d .dmaMHc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.jR8x9d .dmaMHc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before,.jR8x9d .dmaMHc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.jR8x9d .dmaMHc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .dmaMHc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.jR8x9d .dmaMHc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}.jR8x9d .dmaMHc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS{color:rgb(154,160,166)}.jR8x9d .dmaMHc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-clz4Ic{border-bottom-color:rgba(232,234,237,.12)}.jR8x9d .dmaMHc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc{color:rgb(232,234,237)}.jR8x9d .dmaMHc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-pZXsl::before,.jR8x9d .dmaMHc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b .VfPpkd-StrnGf-rymPhb-pZXsl::after{background-color:rgb(232,234,237);background-color:var(--mdc-ripple-color,rgb(232,234,237))}.jR8x9d .dmaMHc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before,.jR8x9d .dmaMHc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.jR8x9d .dmaMHc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before,.jR8x9d .dmaMHc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.jR8x9d .dmaMHc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .dmaMHc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.jR8x9d .dmaMHc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}}@media screen and (prefers-color-scheme:dark) and (-ms-high-contrast:active),screen and (prefers-color-scheme:dark) and (forced-colors:active){.jR8x9d .dmaMHc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c,.jR8x9d .dmaMHc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-fpDzbe-fmcmS,.jR8x9d .dmaMHc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS{color:GrayText}.jR8x9d .dmaMHc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-StrnGf-rymPhb-b9t22c{opacity:1}}@media screen and (prefers-color-scheme:dark){.jR8x9d .dmaMHc .VfPpkd-BFbNVe-bF1uUb{opacity:.08}.jR8x9d .dmaMHc .VfPpkd-rymPhb-Gtdoyb,.jR8x9d .dmaMHc .VfPpkd-rymPhb-fpDzbe-fmcmS{color:rgb(232,234,237)}.jR8x9d .dmaMHc .VfPpkd-rymPhb-L8ivfd-fmcmS,.jR8x9d .dmaMHc .VfPpkd-rymPhb-bC5pod-fmcmS,.jR8x9d .dmaMHc .VfPpkd-rymPhb-JMEf7e{color:rgb(154,160,166)}.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb,.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e,.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-Gtdoyb,.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-fpDzbe-fmcmS,.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-L8ivfd-fmcmS,.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-bC5pod-fmcmS,.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb,.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e,.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e{color:rgb(232,234,237)}.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-KkROqb,.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-Gtdoyb,.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-JMEf7e{opacity:.38}.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-Gtdoyb,.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-fpDzbe-fmcmS,.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-rymPhb-Gtdoyb,.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b .VfPpkd-rymPhb-fpDzbe-fmcmS,.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb,.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b-OWXEXe-pXU01b.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb{color:rgb(232,234,237)}.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::before{opacity:0}.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd{background-color:rgba(138,180,248,.24)}.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::before,.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::after{background-color:rgb(138,180,248);background-color:var(--mdc-ripple-color,rgb(138,180,248))}.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-rymPhb-pZXsl::before,.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-rymPhb-pZXsl::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-rymPhb-pZXsl::before,.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-rymPhb-pZXsl::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-rymPhb-pZXsl::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-rymPhb-pZXsl::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}.jR8x9d .dmaMHc .VfPpkd-rymPhb-L8ivfd-fmcmS{color:rgb(154,160,166)}.jR8x9d .dmaMHc .VfPpkd-rymPhb-clz4Ic{background-color:rgba(232,234,237,.12)}.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb,.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e{color:rgb(232,234,237)}.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::before,.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b .VfPpkd-rymPhb-pZXsl::after{background-color:rgb(232,234,237);background-color:var(--mdc-ripple-color,rgb(232,234,237))}.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b:hover .VfPpkd-rymPhb-pZXsl::before,.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-rymPhb-pZXsl::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-rymPhb-pZXsl::before,.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-rymPhb-pZXsl::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-rymPhb-pZXsl::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-rymPhb-pZXsl::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}}@media screen and (prefers-color-scheme:dark) and (forced-colors:active){.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-Gtdoyb,.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-fpDzbe-fmcmS,.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-L8ivfd-fmcmS,.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-bC5pod-fmcmS,.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb,.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e,.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me.VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-r4m2rf .VfPpkd-rymPhb-JMEf7e{color:GrayText}.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-KkROqb,.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-Gtdoyb,.jR8x9d .dmaMHc .VfPpkd-rymPhb-ibnC6b-OWXEXe-OWB6Me .VfPpkd-rymPhb-JMEf7e{opacity:1}}@media screen and (prefers-color-scheme:dark){.jR8x9d .dmaMHc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-L8ivfd-fmcmS{color:rgb(154,160,166)}.jR8x9d .dmaMHc .VfPpkd-StrnGf-rymPhb .VfPpkd-StrnGf-rymPhb-f7MjDc,.jR8x9d .dmaMHc .VfPpkd-rymPhb .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-M1Soyc-Bz112c .VfPpkd-rymPhb-KkROqb,.jR8x9d .dmaMHc .VfPpkd-rymPhb .VfPpkd-rymPhb-ibnC6b-OWXEXe-SfQLQb-UbuQg-Bz112c .VfPpkd-rymPhb-JMEf7e{color:rgb(232,234,237)}.jR8x9d .dmaMHc .VfPpkd-rymPhb-fpDzbe-fmcmS{letter-spacing:.00625em}.jR8x9d .dmaMHc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd,.jR8x9d .dmaMHc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd{background-color:rgba(242,139,130,.24)}.jR8x9d .dmaMHc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before,.jR8x9d .dmaMHc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::after,.jR8x9d .dmaMHc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::before,.jR8x9d .dmaMHc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-StrnGf-rymPhb-pZXsl::after{background-color:rgb(242,139,130);background-color:var(--mdc-ripple-color,rgb(242,139,130))}.jR8x9d .dmaMHc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before,.jR8x9d .dmaMHc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before,.jR8x9d .dmaMHc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-StrnGf-rymPhb-pZXsl::before,.jR8x9d .dmaMHc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-StrnGf-rymPhb-pZXsl::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.jR8x9d .dmaMHc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before,.jR8x9d .dmaMHc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before,.jR8x9d .dmaMHc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-StrnGf-rymPhb-pZXsl::before,.jR8x9d .dmaMHc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-StrnGf-rymPhb-pZXsl::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.jR8x9d .dmaMHc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after,.jR8x9d .dmaMHc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-StrnGf-rymPhb-pZXsl::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .dmaMHc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after,.jR8x9d .dmaMHc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-StrnGf-rymPhb-pZXsl::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.jR8x9d .dmaMHc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::before,.jR8x9d .dmaMHc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::after,.jR8x9d .dmaMHc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::before,.jR8x9d .dmaMHc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd .VfPpkd-rymPhb-pZXsl::after{background-color:rgb(242,139,130);background-color:var(--mdc-ripple-color,rgb(242,139,130))}.jR8x9d .dmaMHc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-rymPhb-pZXsl::before,.jR8x9d .dmaMHc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-rymPhb-pZXsl::before,.jR8x9d .dmaMHc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:hover .VfPpkd-rymPhb-pZXsl::before,.jR8x9d .dmaMHc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-rymPhb-pZXsl::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.jR8x9d .dmaMHc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-rymPhb-pZXsl::before,.jR8x9d .dmaMHc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-rymPhb-pZXsl::before,.jR8x9d .dmaMHc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-rymPhb-pZXsl::before,.jR8x9d .dmaMHc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-rymPhb-pZXsl::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.jR8x9d .dmaMHc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-rymPhb-pZXsl::after,.jR8x9d .dmaMHc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-rymPhb-pZXsl::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .dmaMHc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-rymPhb-pZXsl::after,.jR8x9d .dmaMHc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-rymPhb-pZXsl::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.jR8x9d .dmaMHc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-StrnGf-rymPhb-ibnC6b.VfPpkd-StrnGf-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d,.jR8x9d .dmaMHc.VfPpkd-YPmvEd-OWXEXe-UJflGc .VfPpkd-rymPhb-ibnC6b.VfPpkd-rymPhb-ibnC6b-OWXEXe-gk6SMd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}.jR8x9d .RnXJS:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-TkwUic{background-color:rgb(60,64,67)}.jR8x9d .RnXJS.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-TkwUic{background-color:rgba(232,234,237,.04)}.jR8x9d .RnXJS:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgb(154,160,166)}.jR8x9d .RnXJS:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):hover .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgb(248,249,250)}.jR8x9d .RnXJS:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::after{border-bottom-color:rgb(138,180,248)}.jR8x9d .RnXJS.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgba(232,234,237,.38)}.jR8x9d .RnXJS:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(189,193,198)}.jR8x9d .RnXJS:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc{color:rgb(138,180,248)}.jR8x9d .RnXJS:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):not(.VfPpkd-O1htCb-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc{color:rgb(248,249,250)}.jR8x9d .RnXJS.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-NLUYnc-V67aGc{color:rgba(232,234,237,.38)}.jR8x9d .RnXJS:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me)+.VfPpkd-O1htCb-W0vJo-fmcmS{color:rgb(154,160,166)}.jR8x9d .RnXJS.VfPpkd-O1htCb-OWXEXe-OWB6Me+.VfPpkd-O1htCb-W0vJo-fmcmS{color:rgba(232,234,237,.38)}.jR8x9d .RnXJS:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-UJflGc+.VfPpkd-O1htCb-W0vJo-fmcmS-OWXEXe-Rfh2Tc-EglORb{color:rgb(246,174,169)}.jR8x9d .RnXJS:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):not(.VfPpkd-O1htCb-OWXEXe-XpnDCe):hover.VfPpkd-O1htCb-OWXEXe-UJflGc+.VfPpkd-O1htCb-W0vJo-fmcmS-OWXEXe-Rfh2Tc-EglORb{color:rgb(246,174,169)}.jR8x9d .RnXJS:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-uusGie-fmcmS{color:rgb(232,234,237)}.jR8x9d .RnXJS.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-uusGie-fmcmS{color:rgba(232,234,237,.38)}}@media screen and (prefers-color-scheme:dark) and (forced-colors:active){.jR8x9d .RnXJS.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-NLUYnc-V67aGc,.jR8x9d .RnXJS.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-uusGie-fmcmS{color:GrayText}}@media screen and (prefers-color-scheme:dark){.jR8x9d .RnXJS:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-t08AT-Bz112c{fill:rgb(189,193,198)}.jR8x9d .RnXJS:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):not(.VfPpkd-O1htCb-OWXEXe-XpnDCe):hover .VfPpkd-t08AT-Bz112c{fill:rgb(248,249,250)}.jR8x9d .RnXJS:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-t08AT-Bz112c{fill:rgb(138,180,248)}.jR8x9d .RnXJS.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-t08AT-Bz112c{fill:rgba(232,234,237,.38)}.jR8x9d .RnXJS:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-cTi5dd{color:rgb(189,193,198)}.jR8x9d .RnXJS.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-cTi5dd{color:rgba(232,234,237,.38)}.jR8x9d .RnXJS.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgb(246,174,169)}.jR8x9d .RnXJS.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):hover .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgb(246,174,169)}.jR8x9d .RnXJS.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::after{border-bottom-color:rgb(246,174,169)}.jR8x9d .RnXJS.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(246,174,169)}.jR8x9d .RnXJS.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):not(.VfPpkd-O1htCb-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc{color:rgb(246,174,169)}.jR8x9d .RnXJS.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{color:rgb(246,174,169)}.jR8x9d .RnXJS.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):not(.VfPpkd-O1htCb-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{color:rgb(246,174,169)}.jR8x9d .RnXJS.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-t08AT-Bz112c{fill:rgb(242,139,130)}.jR8x9d .RnXJS.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):not(.VfPpkd-O1htCb-OWXEXe-XpnDCe):hover .VfPpkd-t08AT-Bz112c{fill:rgb(246,174,169)}.jR8x9d .RnXJS.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-t08AT-Bz112c{fill:rgb(242,139,130)}.jR8x9d .RnXJS .VfPpkd-TkwUic .VfPpkd-woaZLe::before,.jR8x9d .RnXJS .VfPpkd-TkwUic .VfPpkd-woaZLe::after{background-color:rgb(241,243,244);background-color:var(--mdc-ripple-color,rgb(241,243,244))}.jR8x9d .RnXJS .VfPpkd-TkwUic:hover .VfPpkd-woaZLe::before,.jR8x9d .RnXJS .VfPpkd-TkwUic.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-woaZLe::before{opacity:.08;opacity:var(--mdc-ripple-hover-opacity,.08)}.jR8x9d .RnXJS .VfPpkd-TkwUic.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-woaZLe::before,.jR8x9d .RnXJS .VfPpkd-TkwUic:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-woaZLe::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.jR8x9d .RnXJS .VfPpkd-TkwUic:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-woaZLe::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .RnXJS .VfPpkd-TkwUic:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-woaZLe::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.jR8x9d .RnXJS .VfPpkd-TkwUic.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}.jR8x9d .UAQDDf:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Brv4Fb,.jR8x9d .UAQDDf:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Ra9xwd,.jR8x9d .UAQDDf:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-MpmGFe{border-color:rgb(189,193,198)}.jR8x9d .UAQDDf:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):not(.VfPpkd-O1htCb-OWXEXe-XpnDCe) .VfPpkd-TkwUic:hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Brv4Fb,.jR8x9d .UAQDDf:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):not(.VfPpkd-O1htCb-OWXEXe-XpnDCe) .VfPpkd-TkwUic:hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Ra9xwd,.jR8x9d .UAQDDf:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):not(.VfPpkd-O1htCb-OWXEXe-XpnDCe) .VfPpkd-TkwUic:hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-MpmGFe{border-color:rgb(248,249,250)}.jR8x9d .UAQDDf:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Brv4Fb,.jR8x9d .UAQDDf:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Ra9xwd,.jR8x9d .UAQDDf:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-MpmGFe{border-color:rgb(138,180,248)}.jR8x9d .UAQDDf.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-NSFCdd-Brv4Fb,.jR8x9d .UAQDDf.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-NSFCdd-Ra9xwd,.jR8x9d .UAQDDf.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-NSFCdd-MpmGFe{border-color:rgba(232,234,237,.12)}.jR8x9d .UAQDDf:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(154,160,166)}.jR8x9d .UAQDDf:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc{color:rgb(138,180,248)}.jR8x9d .UAQDDf:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):not(.VfPpkd-O1htCb-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc{color:rgb(248,249,250)}.jR8x9d .UAQDDf.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-NLUYnc-V67aGc{color:rgba(232,234,237,.38)}.jR8x9d .UAQDDf:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me)+.VfPpkd-O1htCb-W0vJo-fmcmS{color:rgb(154,160,166)}.jR8x9d .UAQDDf.VfPpkd-O1htCb-OWXEXe-OWB6Me+.VfPpkd-O1htCb-W0vJo-fmcmS{color:rgba(232,234,237,.38)}.jR8x9d .UAQDDf:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-UJflGc+.VfPpkd-O1htCb-W0vJo-fmcmS-OWXEXe-Rfh2Tc-EglORb{color:rgb(242,139,130)}.jR8x9d .UAQDDf:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):not(.VfPpkd-O1htCb-OWXEXe-XpnDCe):hover.VfPpkd-O1htCb-OWXEXe-UJflGc+.VfPpkd-O1htCb-W0vJo-fmcmS-OWXEXe-Rfh2Tc-EglORb{color:rgb(246,174,169)}.jR8x9d .UAQDDf:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-uusGie-fmcmS{color:rgb(232,234,237)}.jR8x9d .UAQDDf.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-uusGie-fmcmS{color:rgba(232,234,237,.38)}}@media screen and (prefers-color-scheme:dark) and (forced-colors:active){.jR8x9d .UAQDDf.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-NLUYnc-V67aGc,.jR8x9d .UAQDDf.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-uusGie-fmcmS{color:GrayText}}@media screen and (prefers-color-scheme:dark){.jR8x9d .UAQDDf:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-t08AT-Bz112c{fill:rgb(154,160,166)}.jR8x9d .UAQDDf:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):not(.VfPpkd-O1htCb-OWXEXe-XpnDCe):hover .VfPpkd-t08AT-Bz112c{fill:rgb(248,249,250)}.jR8x9d .UAQDDf:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-t08AT-Bz112c{fill:rgb(138,180,248)}.jR8x9d .UAQDDf.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-t08AT-Bz112c{fill:rgba(232,234,237,.38)}.jR8x9d .UAQDDf:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-cTi5dd{color:rgb(154,160,166)}.jR8x9d .UAQDDf.VfPpkd-O1htCb-OWXEXe-OWB6Me .VfPpkd-cTi5dd{color:rgba(232,234,237,.38)}.jR8x9d .UAQDDf.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Brv4Fb,.jR8x9d .UAQDDf.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Ra9xwd,.jR8x9d .UAQDDf.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-MpmGFe{border-color:rgb(242,139,130)}.jR8x9d .UAQDDf.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):not(.VfPpkd-O1htCb-OWXEXe-XpnDCe) .VfPpkd-TkwUic:hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Brv4Fb,.jR8x9d .UAQDDf.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):not(.VfPpkd-O1htCb-OWXEXe-XpnDCe) .VfPpkd-TkwUic:hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Ra9xwd,.jR8x9d .UAQDDf.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):not(.VfPpkd-O1htCb-OWXEXe-XpnDCe) .VfPpkd-TkwUic:hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-MpmGFe{border-color:rgb(246,174,169)}.jR8x9d .UAQDDf.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Brv4Fb,.jR8x9d .UAQDDf.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Ra9xwd,.jR8x9d .UAQDDf.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-MpmGFe{border-color:rgb(242,139,130)}.jR8x9d .UAQDDf.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(242,139,130)}.jR8x9d .UAQDDf.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):not(.VfPpkd-O1htCb-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc{color:rgb(246,174,169)}.jR8x9d .UAQDDf.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{color:rgb(242,139,130)}.jR8x9d .UAQDDf.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):not(.VfPpkd-O1htCb-OWXEXe-XpnDCe):hover .VfPpkd-NLUYnc-V67aGc-OWXEXe-TATcMc-KLRBe{color:rgb(246,174,169)}.jR8x9d .UAQDDf.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me) .VfPpkd-t08AT-Bz112c{fill:rgb(242,139,130)}.jR8x9d .UAQDDf.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me):not(.VfPpkd-O1htCb-OWXEXe-XpnDCe):hover .VfPpkd-t08AT-Bz112c{fill:rgb(246,174,169)}.jR8x9d .UAQDDf.VfPpkd-O1htCb-OWXEXe-UJflGc:not(.VfPpkd-O1htCb-OWXEXe-OWB6Me).VfPpkd-O1htCb-OWXEXe-XpnDCe .VfPpkd-t08AT-Bz112c{fill:rgb(242,139,130)}.jR8x9d .UlwoYd .VfPpkd-UTM9ec-tmWYNe{background-color:rgb(138,180,248);border-color:rgb(138,180,248)}.jR8x9d .UlwoYd .VfPpkd-UTM9ec-OWXEXe-ma6Yeb .VfPpkd-UTM9ec-tmWYNe,.jR8x9d .UlwoYd .VfPpkd-UTM9ec-OWXEXe-ma6Yeb.VfPpkd-UTM9ec:hover .VfPpkd-UTM9ec-tmWYNe,.jR8x9d .UlwoYd .VfPpkd-UTM9ec-OWXEXe-ma6Yeb.VfPpkd-UTM9ec-OWXEXe-XpnDCe .VfPpkd-UTM9ec-tmWYNe{border-color:#fff}.jR8x9d .UlwoYd.VfPpkd-SxecR-OWXEXe-OWB6Me .VfPpkd-UTM9ec-tmWYNe{background-color:rgb(232,234,237);border-color:rgb(232,234,237)}.jR8x9d .UlwoYd.VfPpkd-SxecR-OWXEXe-OWB6Me .VfPpkd-UTM9ec-OWXEXe-ma6Yeb .VfPpkd-UTM9ec-tmWYNe,.jR8x9d .UlwoYd.VfPpkd-SxecR-OWXEXe-OWB6Me .VfPpkd-UTM9ec-OWXEXe-ma6Yeb.VfPpkd-UTM9ec:hover .VfPpkd-UTM9ec-tmWYNe,.jR8x9d .UlwoYd.VfPpkd-SxecR-OWXEXe-OWB6Me .VfPpkd-UTM9ec-OWXEXe-ma6Yeb.VfPpkd-UTM9ec-OWXEXe-XpnDCe .VfPpkd-UTM9ec-tmWYNe{border-color:#fff}.jR8x9d .UlwoYd .VfPpkd-UTM9ec::before,.jR8x9d .UlwoYd .VfPpkd-UTM9ec::after{background-color:rgb(138,180,248);background-color:var(--mdc-ripple-color,rgb(138,180,248))}.jR8x9d .UlwoYd .VfPpkd-UTM9ec:hover::before,.jR8x9d .UlwoYd .VfPpkd-UTM9ec.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE::before{opacity:.08;opacity:var(--mdc-ripple-hover-opacity,.08)}.jR8x9d .UlwoYd .VfPpkd-UTM9ec.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe::before,.jR8x9d .UlwoYd .VfPpkd-UTM9ec:not(.VfPpkd-ksKsZd-mWPk3d):focus::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.24;opacity:var(--mdc-ripple-focus-opacity,.24)}.jR8x9d .UlwoYd .VfPpkd-UTM9ec:not(.VfPpkd-ksKsZd-mWPk3d)::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .UlwoYd .VfPpkd-UTM9ec:not(.VfPpkd-ksKsZd-mWPk3d):active::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.24;opacity:var(--mdc-ripple-press-opacity,.24)}.jR8x9d .UlwoYd .VfPpkd-UTM9ec.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.24)}.jR8x9d .UlwoYd .VfPpkd-UTM9ec:hover .VfPpkd-UTM9ec-tmWYNe,.jR8x9d .UlwoYd .VfPpkd-UTM9ec-OWXEXe-XpnDCe .VfPpkd-UTM9ec-tmWYNe{background-color:rgb(210,227,252);border-color:rgb(210,227,252)}.jR8x9d .UlwoYd .VfPpkd-UTM9ec:hover .VfPpkd-UTM9ec-OWXEXe-ma6Yeb .VfPpkd-UTM9ec-tmWYNe,.jR8x9d .UlwoYd .VfPpkd-UTM9ec:hover .VfPpkd-UTM9ec-OWXEXe-ma6Yeb.VfPpkd-UTM9ec:hover .VfPpkd-UTM9ec-tmWYNe,.jR8x9d .UlwoYd .VfPpkd-UTM9ec:hover .VfPpkd-UTM9ec-OWXEXe-ma6Yeb.VfPpkd-UTM9ec-OWXEXe-XpnDCe .VfPpkd-UTM9ec-tmWYNe,.jR8x9d .UlwoYd .VfPpkd-UTM9ec-OWXEXe-XpnDCe .VfPpkd-UTM9ec-OWXEXe-ma6Yeb .VfPpkd-UTM9ec-tmWYNe,.jR8x9d .UlwoYd .VfPpkd-UTM9ec-OWXEXe-XpnDCe .VfPpkd-UTM9ec-OWXEXe-ma6Yeb.VfPpkd-UTM9ec:hover .VfPpkd-UTM9ec-tmWYNe,.jR8x9d .UlwoYd .VfPpkd-UTM9ec-OWXEXe-XpnDCe .VfPpkd-UTM9ec-OWXEXe-ma6Yeb.VfPpkd-UTM9ec-OWXEXe-XpnDCe .VfPpkd-UTM9ec-tmWYNe{border-color:#fff}.jR8x9d .UlwoYd .VfPpkd-yCQwvc-OWXEXe-bp49T{border-color:rgb(138,180,248)}.jR8x9d .UlwoYd.VfPpkd-SxecR-OWXEXe-OWB6Me .VfPpkd-yCQwvc-OWXEXe-bp49T{border-color:rgb(232,234,237)}.jR8x9d .UlwoYd .VfPpkd-yCQwvc-OWXEXe-mt1Mkb{background-color:rgb(32,33,36);opacity:1}.jR8x9d .UlwoYd.VfPpkd-SxecR-OWXEXe-OWB6Me .VfPpkd-yCQwvc-OWXEXe-mt1Mkb{background-color:rgba(232,234,237,.38);opacity:1}.jR8x9d .UlwoYd .VfPpkd-zD2WHb-SYOSDb-OWXEXe-auswjd,.jR8x9d .UlwoYd.VfPpkd-SxecR-OWXEXe-OWB6Me .VfPpkd-zD2WHb-SYOSDb-OWXEXe-auswjd{background-color:rgb(32,33,36);opacity:.38}}@media screen and (prefers-color-scheme:dark) and (forced-colors:active){.jR8x9d .UlwoYd .VfPpkd-zD2WHb-SYOSDb-OWXEXe-auswjd{background-color:Canvas;opacity:1}}@media screen and (prefers-color-scheme:dark){.jR8x9d .UlwoYd .VfPpkd-zD2WHb-SYOSDb-OWXEXe-mt1Mkb{background-color:rgb(138,180,248);opacity:.38}.jR8x9d .UlwoYd.VfPpkd-SxecR-OWXEXe-OWB6Me .VfPpkd-zD2WHb-SYOSDb-OWXEXe-mt1Mkb{background-color:rgb(232,234,237);opacity:.38}}@media screen and (prefers-color-scheme:dark) and (forced-colors:active){.jR8x9d .UlwoYd .VfPpkd-zD2WHb-SYOSDb-OWXEXe-mt1Mkb{background-color:CanvasText;opacity:1}}@media screen and (prefers-color-scheme:dark){.jR8x9d .UlwoYd:not(.VfPpkd-SxecR-OWXEXe-OWB6Me) .VfPpkd-yCQwvc-OWXEXe-mt1Mkb::before{background-color:rgba(138,180,248,.24);border-radius:inherit;content:"";height:100%;position:absolute;width:100%}.jR8x9d .UlwoYd .VfPpkd-MIfjnf-uDEFge{background-color:rgb(138,180,248);opacity:1}.jR8x9d .UlwoYd .VfPpkd-MIfjnf-uDEFge::before{border-top-color:rgb(138,180,248)}.jR8x9d .UlwoYd .VfPpkd-MIfjnf-uDEFge{color:rgb(32,33,36)}.jR8x9d .UlwoYd.VfPpkd-SxecR .VfPpkd-yCQwvc-OWXEXe-bp49T{-webkit-transform-origin:left;transform-origin:left}.jR8x9d .UlwoYd .VfPpkd-MIfjnf-uDEFge{border-radius:16px;height:28px;padding:0 8px}.jR8x9d .UlwoYd .VfPpkd-MIfjnf-uDEFge-fmcmS{font-family:"Roboto Mono",Roboto,sans-serif;font-size:.75rem;font-weight:500;white-space:nowrap}.jR8x9d .UlwoYd .VfPpkd-UTM9ec.VfPpkd-UTM9ec-OWXEXe-fmcmS-YuD1xf-lTBxed .VfPpkd-MIfjnf-uDEFge-fmcmS{font-family:Roboto,sans-serif}.jR8x9d .UlwoYd .VfPpkd-UTM9ec.VfPpkd-UTM9ec-OWXEXe-Wetbn-lTBxed .VfPpkd-MIfjnf-uDEFge-haAclf{bottom:40px;-webkit-transform:rotate(-45deg);transform:rotate(-45deg);-webkit-transform-origin:bottom left;transform-origin:bottom left}.jR8x9d .UlwoYd .VfPpkd-UTM9ec.VfPpkd-UTM9ec-OWXEXe-Wetbn-lTBxed .VfPpkd-MIfjnf-uDEFge{border-radius:50% 50% 50% 0;height:28px;-webkit-box-pack:center;-webkit-justify-content:center;justify-content:center;padding:0;position:relative;width:28px}.jR8x9d .UlwoYd .VfPpkd-UTM9ec.VfPpkd-UTM9ec-OWXEXe-Wetbn-lTBxed .VfPpkd-MIfjnf-uDEFge::before{display:none}.jR8x9d .UlwoYd .VfPpkd-UTM9ec.VfPpkd-UTM9ec-OWXEXe-Wetbn-lTBxed .VfPpkd-MIfjnf-uDEFge-fmcmS{-webkit-transform:rotate(45deg);transform:rotate(45deg)}.jR8x9d .TFhMef .VfPpkd-YAxtVc{background-color:#fff}.jR8x9d .TFhMef .VfPpkd-gIZMF{color:rgb(60,64,67)}.jR8x9d .TFhMef .VfPpkd-IkaYrd:not(:disabled){background-color:transparent}.jR8x9d .TFhMef .VfPpkd-IkaYrd:not(:disabled){color:rgb(26,115,232);color:var(--gm-colortextbutton-ink-color,rgb(26,115,232))}.jR8x9d .TFhMef .VfPpkd-IkaYrd:disabled{color:rgba(60,64,67,.38);color:var(--gm-colortextbutton-disabled-ink-color,rgba(60,64,67,.38))}.jR8x9d .TFhMef .VfPpkd-IkaYrd .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo,.jR8x9d .TFhMef .VfPpkd-IkaYrd .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:rgb(26,115,232)}}@media screen and (prefers-color-scheme:dark) and (-ms-high-contrast:active),screen and (prefers-color-scheme:dark) and (forced-colors:active){.jR8x9d .TFhMef .VfPpkd-IkaYrd .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-uI4vCe-LkdAo,.jR8x9d .TFhMef .VfPpkd-IkaYrd .VfPpkd-UdE5de-uDEFge .VfPpkd-JGcpL-IdXvz-LkdAo-Bd00G{stroke:CanvasText}}@media screen and (prefers-color-scheme:dark){.jR8x9d .TFhMef .VfPpkd-IkaYrd:hover:not(:disabled),.jR8x9d .TFhMef .VfPpkd-IkaYrd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:disabled),.jR8x9d .TFhMef .VfPpkd-IkaYrd:not(.VfPpkd-ksKsZd-mWPk3d):focus:not(:disabled),.jR8x9d .TFhMef .VfPpkd-IkaYrd:active:not(:disabled){color:rgb(23,78,166);color:var(--gm-colortextbutton-ink-color--stateful,rgb(23,78,166))}.jR8x9d .TFhMef .VfPpkd-IkaYrd .VfPpkd-Jh9lGc::before,.jR8x9d .TFhMef .VfPpkd-IkaYrd .VfPpkd-Jh9lGc::after{background-color:rgb(26,115,232);background-color:var(--gm-colortextbutton-state-color,rgb(26,115,232))}.jR8x9d .TFhMef .VfPpkd-IkaYrd:hover .VfPpkd-Jh9lGc::before,.jR8x9d .TFhMef .VfPpkd-IkaYrd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.jR8x9d .TFhMef .VfPpkd-IkaYrd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.jR8x9d .TFhMef .VfPpkd-IkaYrd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.jR8x9d .TFhMef .VfPpkd-IkaYrd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .TFhMef .VfPpkd-IkaYrd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-press-opacity,.12)}.jR8x9d .TFhMef .VfPpkd-IkaYrd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.12)}.jR8x9d .TFhMef .VfPpkd-IkaYrd:disabled:hover .VfPpkd-Jh9lGc::before,.jR8x9d .TFhMef .VfPpkd-IkaYrd:disabled.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Jh9lGc::before{opacity:0;opacity:var(--mdc-ripple-hover-opacity,0)}.jR8x9d .TFhMef .VfPpkd-IkaYrd:disabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Jh9lGc::before,.jR8x9d .TFhMef .VfPpkd-IkaYrd:disabled:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:0;opacity:var(--mdc-ripple-focus-opacity,0)}.jR8x9d .TFhMef .VfPpkd-IkaYrd:disabled:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .TFhMef .VfPpkd-IkaYrd:disabled:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:0;opacity:var(--mdc-ripple-press-opacity,0)}.jR8x9d .TFhMef .VfPpkd-IkaYrd:disabled.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0)}.jR8x9d .TFhMef .VfPpkd-TolmDb{color:rgb(60,64,67);z-index:0}.jR8x9d .TFhMef .VfPpkd-TolmDb .VfPpkd-Bz112c-Jh9lGc::before,.jR8x9d .TFhMef .VfPpkd-TolmDb .VfPpkd-Bz112c-Jh9lGc::after{background-color:rgb(60,64,67);background-color:var(--mdc-ripple-color,rgb(60,64,67))}.jR8x9d .TFhMef .VfPpkd-TolmDb:hover .VfPpkd-Bz112c-Jh9lGc::before,.jR8x9d .TFhMef .VfPpkd-TolmDb.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Bz112c-Jh9lGc::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.jR8x9d .TFhMef .VfPpkd-TolmDb.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Bz112c-Jh9lGc::before,.jR8x9d .TFhMef .VfPpkd-TolmDb:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Bz112c-Jh9lGc::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.jR8x9d .TFhMef .VfPpkd-TolmDb:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Bz112c-Jh9lGc::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .TFhMef .VfPpkd-TolmDb:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Bz112c-Jh9lGc::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-press-opacity,.12)}.jR8x9d .TFhMef .VfPpkd-TolmDb.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.12)}.jR8x9d .TFhMef .VfPpkd-TolmDb .VfPpkd-Bz112c-Jh9lGc::before,.jR8x9d .TFhMef .VfPpkd-TolmDb .VfPpkd-Bz112c-Jh9lGc::after{z-index:-1}.jR8x9d .TFhMef .VfPpkd-TolmDb:disabled{color:rgba(60,64,67,.38);color:var(--gm-iconbutton-disabled-ink-color,rgba(60,64,67,.38))}.jR8x9d .pBHsAc{width:36px}.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled .VfPpkd-uMhiad::after{background:rgb(138,180,248)}.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe):not(:active) .VfPpkd-uMhiad::after{background:rgb(174,203,250)}.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:active) .VfPpkd-uMhiad::after{background:rgb(174,203,250)}.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:active .VfPpkd-uMhiad::after{background:rgb(174,203,250)}.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-gk6SMd:disabled .VfPpkd-uMhiad::after{background:rgb(232,234,237)}.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-uqeOfd:enabled .VfPpkd-uMhiad::after{background:rgb(154,160,166)}.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-uqeOfd:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe):not(:active) .VfPpkd-uMhiad::after{background:rgb(248,249,250)}.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-uqeOfd:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:active) .VfPpkd-uMhiad::after{background:rgb(248,249,250)}.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-uqeOfd:enabled:active .VfPpkd-uMhiad::after{background:rgb(248,249,250)}.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-uqeOfd:disabled .VfPpkd-uMhiad::after{background:rgb(232,234,237)}.jR8x9d .pBHsAc .VfPpkd-uMhiad::before{background:rgb(32,33,36)}.jR8x9d .pBHsAc:enabled .VfPpkd-VRSVNe{box-shadow:0 1px 2px 0 rgba(0,0,0,.3),0 1px 3px 1px rgba(0,0,0,.15)}.jR8x9d .pBHsAc:enabled .VfPpkd-VRSVNe .VfPpkd-BFbNVe-bF1uUb{opacity:.05}.jR8x9d .pBHsAc:enabled .VfPpkd-VRSVNe .VfPpkd-BFbNVe-bF1uUb{background-color:rgb(232,234,237)}.jR8x9d .pBHsAc:disabled .VfPpkd-VRSVNe{box-shadow:none}.jR8x9d .pBHsAc:disabled .VfPpkd-VRSVNe .VfPpkd-BFbNVe-bF1uUb{opacity:0}.jR8x9d .pBHsAc:disabled .VfPpkd-VRSVNe .VfPpkd-BFbNVe-bF1uUb{background-color:rgb(232,234,237)}.jR8x9d .pBHsAc .VfPpkd-DVBDLb-LhBDec-sM5MNb,.jR8x9d .pBHsAc .VfPpkd-uMhiad{height:20px}.jR8x9d .pBHsAc:disabled .VfPpkd-uMhiad::after{opacity:.38}.jR8x9d .pBHsAc .VfPpkd-uMhiad{border-radius:10px 10px 10px 10px}.jR8x9d .pBHsAc .VfPpkd-uMhiad{width:20px}.jR8x9d .pBHsAc .VfPpkd-uMhiad-u014N{width:calc(100% - 20px)}.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled .VfPpkd-pafCAf{fill:rgb(32,33,36)}.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-gk6SMd:disabled .VfPpkd-pafCAf{fill:rgb(32,33,36)}.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-uqeOfd:enabled .VfPpkd-pafCAf{fill:rgb(32,33,36)}.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-uqeOfd:disabled .VfPpkd-pafCAf{fill:rgb(32,33,36)}.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-gk6SMd:disabled .VfPpkd-lw9akd{opacity:.38}.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-uqeOfd:disabled .VfPpkd-lw9akd{opacity:.38}.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-gk6SMd .VfPpkd-pafCAf,.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-uqeOfd .VfPpkd-pafCAf{width:18px;height:18px}.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe) .VfPpkd-Qsb3yd::before,.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe) .VfPpkd-Qsb3yd::after{background-color:rgb(138,180,248)}.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Qsb3yd::before,.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Qsb3yd::after{background-color:rgb(138,180,248)}.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:active .VfPpkd-Qsb3yd::before,.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:active .VfPpkd-Qsb3yd::after{background-color:rgb(138,180,248)}.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-uqeOfd:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe) .VfPpkd-Qsb3yd::before,.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-uqeOfd:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe) .VfPpkd-Qsb3yd::after{background-color:rgb(232,234,237)}.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-uqeOfd:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Qsb3yd::before,.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-uqeOfd:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Qsb3yd::after{background-color:rgb(232,234,237)}.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-uqeOfd:enabled:active .VfPpkd-Qsb3yd::before,.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-uqeOfd:enabled:active .VfPpkd-Qsb3yd::after{background-color:rgb(232,234,237)}.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe):hover .VfPpkd-Qsb3yd::before,.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe).VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Qsb3yd::before{opacity:.04}.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Qsb3yd::before,.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Qsb3yd::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12}.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:active:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Qsb3yd::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:active:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Qsb3yd::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1}.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled:active.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-switch-selected-pressed-state-layer-opacity,0.1)}.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-uqeOfd:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe):hover .VfPpkd-Qsb3yd::before,.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-uqeOfd:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe).VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-Qsb3yd::before{opacity:.04}.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-uqeOfd:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-Qsb3yd::before,.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-uqeOfd:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-Qsb3yd::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12}.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-uqeOfd:enabled:active:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-Qsb3yd::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-uqeOfd:enabled:active:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-Qsb3yd::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1}.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-uqeOfd:enabled:active.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-switch-unselected-pressed-state-layer-opacity,0.1)}.jR8x9d .pBHsAc .VfPpkd-Qsb3yd{height:48px;width:48px}.jR8x9d .pBHsAc .VfPpkd-l6JLsf{height:14px}.jR8x9d .pBHsAc:disabled .VfPpkd-l6JLsf{opacity:.12}.jR8x9d .pBHsAc:enabled .VfPpkd-l6JLsf::after{background:rgb(26,115,232)}.jR8x9d .pBHsAc:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe):not(:active) .VfPpkd-l6JLsf::after{background:rgb(26,115,232)}.jR8x9d .pBHsAc:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:active) .VfPpkd-l6JLsf::after{background:rgb(26,115,232)}.jR8x9d .pBHsAc:enabled:active .VfPpkd-l6JLsf::after{background:rgb(26,115,232)}.jR8x9d .pBHsAc:disabled .VfPpkd-l6JLsf::after{background:rgb(232,234,237)}.jR8x9d .pBHsAc:enabled .VfPpkd-l6JLsf::before{background:rgb(95,99,104)}.jR8x9d .pBHsAc:enabled:hover:not(.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe):not(:active) .VfPpkd-l6JLsf::before{background:rgb(95,99,104)}.jR8x9d .pBHsAc:enabled.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe:not(:active) .VfPpkd-l6JLsf::before{background:rgb(95,99,104)}.jR8x9d .pBHsAc:enabled:active .VfPpkd-l6JLsf::before{background:rgb(95,99,104)}.jR8x9d .pBHsAc:disabled .VfPpkd-l6JLsf::before{background:rgb(232,234,237)}.jR8x9d .pBHsAc .VfPpkd-l6JLsf{border-radius:7px 7px 7px 7px}}@media screen and (prefers-color-scheme:dark) and (-ms-high-contrast:active),screen and (prefers-color-scheme:dark) and (forced-colors:active){.jR8x9d .pBHsAc:disabled .VfPpkd-uMhiad::after{opacity:1}.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-gk6SMd:enabled .VfPpkd-pafCAf{fill:ButtonText}.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-gk6SMd:disabled .VfPpkd-pafCAf{fill:GrayText}.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-uqeOfd:enabled .VfPpkd-pafCAf{fill:ButtonText}.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-uqeOfd:disabled .VfPpkd-pafCAf{fill:GrayText}.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-gk6SMd:disabled .VfPpkd-lw9akd{opacity:1}.jR8x9d .pBHsAc.VfPpkd-scr2fc-OWXEXe-uqeOfd:disabled .VfPpkd-lw9akd{opacity:1}.jR8x9d .pBHsAc:disabled .VfPpkd-l6JLsf{opacity:1}}@media screen and (prefers-color-scheme:dark){.jR8x9d .FEsNhd{font-family:"Google Sans",Roboto,Arial,sans-serif;line-height:1.25rem;font-size:.875rem;letter-spacing:.0178571429em;font-weight:500;padding-right:16px;padding-left:16px;text-transform:none;min-width:auto}.jR8x9d .FEsNhd .VfPpkd-jY41G-V67aGc{color:rgb(154,160,166)}.jR8x9d .FEsNhd .VfPpkd-cfyjzb{color:rgb(154,160,166);fill:currentColor}.jR8x9d .FEsNhd:hover .VfPpkd-YVzG2b::before,.jR8x9d .FEsNhd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-YVzG2b::before{opacity:.08;opacity:var(--mdc-ripple-hover-opacity,.08)}.jR8x9d .FEsNhd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-YVzG2b::before,.jR8x9d .FEsNhd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-YVzG2b::before{opacity:.24;opacity:var(--mdc-ripple-focus-opacity,.24)}.jR8x9d .FEsNhd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-YVzG2b::after{opacity:.24;opacity:var(--mdc-ripple-press-opacity,.24)}.jR8x9d .FEsNhd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.24)}.jR8x9d .FEsNhd:hover .VfPpkd-jY41G-V67aGc,.jR8x9d .FEsNhd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-jY41G-V67aGc,.jR8x9d .FEsNhd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-jY41G-V67aGc,.jR8x9d .FEsNhd:active .VfPpkd-jY41G-V67aGc{color:rgb(232,234,237)}.jR8x9d .FEsNhd:hover .VfPpkd-cfyjzb,.jR8x9d .FEsNhd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-cfyjzb,.jR8x9d .FEsNhd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-cfyjzb,.jR8x9d .FEsNhd:active .VfPpkd-cfyjzb{color:rgb(232,234,237);fill:currentColor}.jR8x9d .FEsNhd .VfPpkd-YVzG2b::before,.jR8x9d .FEsNhd .VfPpkd-YVzG2b::after{background-color:rgb(232,234,237);background-color:var(--mdc-ripple-color,rgb(232,234,237))}.jR8x9d .FEsNhd:hover .VfPpkd-YVzG2b::before,.jR8x9d .FEsNhd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-YVzG2b::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.jR8x9d .FEsNhd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-YVzG2b::before,.jR8x9d .FEsNhd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-YVzG2b::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.jR8x9d .FEsNhd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-YVzG2b::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .FEsNhd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-YVzG2b::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.jR8x9d .FEsNhd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}.jR8x9d .FEsNhd.VfPpkd-AznF2e-OWXEXe-auswjd:hover .VfPpkd-YVzG2b::before,.jR8x9d .FEsNhd.VfPpkd-AznF2e-OWXEXe-auswjd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-YVzG2b::before{opacity:.08;opacity:var(--mdc-ripple-hover-opacity,.08)}.jR8x9d .FEsNhd.VfPpkd-AznF2e-OWXEXe-auswjd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-YVzG2b::before,.jR8x9d .FEsNhd.VfPpkd-AznF2e-OWXEXe-auswjd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-YVzG2b::before{opacity:.24;opacity:var(--mdc-ripple-focus-opacity,.24)}.jR8x9d .FEsNhd.VfPpkd-AznF2e-OWXEXe-auswjd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-YVzG2b::after{opacity:.24;opacity:var(--mdc-ripple-press-opacity,.24)}.jR8x9d .FEsNhd.VfPpkd-AznF2e-OWXEXe-auswjd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.24)}.jR8x9d .FEsNhd.VfPpkd-AznF2e-OWXEXe-auswjd .VfPpkd-jY41G-V67aGc{color:rgb(138,180,248)}.jR8x9d .FEsNhd.VfPpkd-AznF2e-OWXEXe-auswjd .VfPpkd-cfyjzb{color:rgb(138,180,248);fill:currentColor}.jR8x9d .FEsNhd:hover.VfPpkd-AznF2e-OWXEXe-auswjd .VfPpkd-jY41G-V67aGc,.jR8x9d .FEsNhd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-AznF2e-OWXEXe-auswjd .VfPpkd-jY41G-V67aGc,.jR8x9d .FEsNhd:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-AznF2e-OWXEXe-auswjd .VfPpkd-jY41G-V67aGc,.jR8x9d .FEsNhd:active.VfPpkd-AznF2e-OWXEXe-auswjd .VfPpkd-jY41G-V67aGc{color:rgb(174,203,250)}.jR8x9d .FEsNhd:hover.VfPpkd-AznF2e-OWXEXe-auswjd .VfPpkd-cfyjzb,.jR8x9d .FEsNhd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe.VfPpkd-AznF2e-OWXEXe-auswjd .VfPpkd-cfyjzb,.jR8x9d .FEsNhd:not(.VfPpkd-ksKsZd-mWPk3d):focus.VfPpkd-AznF2e-OWXEXe-auswjd .VfPpkd-cfyjzb,.jR8x9d .FEsNhd:active.VfPpkd-AznF2e-OWXEXe-auswjd .VfPpkd-cfyjzb{color:rgb(174,203,250);fill:currentColor}.jR8x9d .FEsNhd:hover .VfPpkd-AznF2e-wEcVzc-OWXEXe-NowJzb,.jR8x9d .FEsNhd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-AznF2e-wEcVzc-OWXEXe-NowJzb,.jR8x9d .FEsNhd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-AznF2e-wEcVzc-OWXEXe-NowJzb,.jR8x9d .FEsNhd:active .VfPpkd-AznF2e-wEcVzc-OWXEXe-NowJzb{border-color:rgb(174,203,250)}.jR8x9d .FEsNhd.VfPpkd-AznF2e-OWXEXe-auswjd .VfPpkd-YVzG2b::before,.jR8x9d .FEsNhd.VfPpkd-AznF2e-OWXEXe-auswjd .VfPpkd-YVzG2b::after{background-color:rgb(174,203,250);background-color:var(--mdc-ripple-color,rgb(174,203,250))}.jR8x9d .FEsNhd.VfPpkd-AznF2e-OWXEXe-auswjd:hover .VfPpkd-YVzG2b::before,.jR8x9d .FEsNhd.VfPpkd-AznF2e-OWXEXe-auswjd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-YVzG2b::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.jR8x9d .FEsNhd.VfPpkd-AznF2e-OWXEXe-auswjd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-YVzG2b::before,.jR8x9d .FEsNhd.VfPpkd-AznF2e-OWXEXe-auswjd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-YVzG2b::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.jR8x9d .FEsNhd.VfPpkd-AznF2e-OWXEXe-auswjd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-YVzG2b::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .FEsNhd.VfPpkd-AznF2e-OWXEXe-auswjd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-YVzG2b::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.jR8x9d .FEsNhd.VfPpkd-AznF2e-OWXEXe-auswjd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}.jR8x9d .V0XHEd{font-family:"Google Sans",Roboto,Arial,sans-serif;line-height:1.25rem;font-size:.875rem;letter-spacing:.0178571429em;font-weight:500;padding-right:16px;padding-left:16px;text-transform:none;min-width:auto}.jR8x9d .V0XHEd .VfPpkd-jY41G-V67aGc{color:rgb(154,160,166)}.jR8x9d .V0XHEd .VfPpkd-cfyjzb{color:rgb(154,160,166);fill:currentColor}.jR8x9d .V0XHEd:hover .VfPpkd-jY41G-V67aGc,.jR8x9d .V0XHEd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-jY41G-V67aGc,.jR8x9d .V0XHEd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-jY41G-V67aGc,.jR8x9d .V0XHEd:active .VfPpkd-jY41G-V67aGc{color:rgb(232,234,237)}.jR8x9d .V0XHEd:hover .VfPpkd-cfyjzb,.jR8x9d .V0XHEd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-cfyjzb,.jR8x9d .V0XHEd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-cfyjzb,.jR8x9d .V0XHEd:active .VfPpkd-cfyjzb{color:rgb(232,234,237);fill:currentColor}.jR8x9d .V0XHEd:hover .VfPpkd-YVzG2b::before,.jR8x9d .V0XHEd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-YVzG2b::before{opacity:.08;opacity:var(--mdc-ripple-hover-opacity,.08)}.jR8x9d .V0XHEd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-YVzG2b::before,.jR8x9d .V0XHEd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-YVzG2b::before{opacity:.24;opacity:var(--mdc-ripple-focus-opacity,.24)}.jR8x9d .V0XHEd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-YVzG2b::after{opacity:.24;opacity:var(--mdc-ripple-press-opacity,.24)}.jR8x9d .V0XHEd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.24)}.jR8x9d .V0XHEd.VfPpkd-AznF2e-OWXEXe-auswjd .VfPpkd-jY41G-V67aGc{color:rgb(232,234,237)}.jR8x9d .V0XHEd.VfPpkd-AznF2e-OWXEXe-auswjd .VfPpkd-cfyjzb{color:rgb(232,234,237);fill:currentColor}.jR8x9d .V0XHEd:hover .VfPpkd-AznF2e-wEcVzc-OWXEXe-NowJzb,.jR8x9d .V0XHEd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-AznF2e-wEcVzc-OWXEXe-NowJzb,.jR8x9d .V0XHEd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-AznF2e-wEcVzc-OWXEXe-NowJzb,.jR8x9d .V0XHEd:active .VfPpkd-AznF2e-wEcVzc-OWXEXe-NowJzb{border-color:rgb(174,203,250)}.jR8x9d .V0XHEd .VfPpkd-YVzG2b::before,.jR8x9d .V0XHEd .VfPpkd-YVzG2b::after{background-color:rgb(232,234,237);background-color:var(--mdc-ripple-color,rgb(232,234,237))}.jR8x9d .V0XHEd:hover .VfPpkd-YVzG2b::before,.jR8x9d .V0XHEd.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-YVzG2b::before{opacity:.04;opacity:var(--mdc-ripple-hover-opacity,.04)}.jR8x9d .V0XHEd.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-YVzG2b::before,.jR8x9d .V0XHEd:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-YVzG2b::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.12;opacity:var(--mdc-ripple-focus-opacity,.12)}.jR8x9d .V0XHEd:not(.VfPpkd-ksKsZd-mWPk3d) .VfPpkd-YVzG2b::after{-webkit-transition:opacity .15s linear;transition:opacity .15s linear}.jR8x9d .V0XHEd:not(.VfPpkd-ksKsZd-mWPk3d):active .VfPpkd-YVzG2b::after{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:.1;opacity:var(--mdc-ripple-press-opacity,.1)}.jR8x9d .V0XHEd.VfPpkd-ksKsZd-mWPk3d{--mdc-ripple-fg-opacity:var(--mdc-ripple-press-opacity,0.1)}.jR8x9d .kte1hc .VfPpkd-AznF2e-wEcVzc-OWXEXe-NowJzb{border-color:rgb(138,180,248)}.jR8x9d .kte1hc .VfPpkd-AznF2e-wEcVzc-OWXEXe-NowJzb{border-top-width:3px}.jR8x9d .kte1hc .VfPpkd-AznF2e-wEcVzc-OWXEXe-NowJzb{border-top-left-radius:3px;border-top-right-radius:3px}.jR8x9d .p4biwf .VfPpkd-AznF2e-wEcVzc-OWXEXe-NowJzb{border-color:rgb(138,180,248)}.jR8x9d .gOPnwc:hover .VfPpkd-fmcmS-OyKIhb::before,.jR8x9d .gOPnwc.VfPpkd-ksKsZd-XxIAqe-OWXEXe-ZmdkE .VfPpkd-fmcmS-OyKIhb::before{opacity:.08;opacity:var(--mdc-ripple-hover-opacity,.08)}.jR8x9d .gOPnwc.VfPpkd-ksKsZd-mWPk3d-OWXEXe-AHe6Kc-XpnDCe .VfPpkd-fmcmS-OyKIhb::before,.jR8x9d .gOPnwc:not(.VfPpkd-ksKsZd-mWPk3d):focus .VfPpkd-fmcmS-OyKIhb::before{-webkit-transition-duration:75ms;transition-duration:75ms;opacity:0;opacity:var(--mdc-ripple-focus-opacity,0)}.jR8x9d .gOPnwc .VfPpkd-fmcmS-OyKIhb::before,.jR8x9d .gOPnwc .VfPpkd-fmcmS-OyKIhb::after{background-color:rgb(241,243,244);background-color:var(--mdc-ripple-color,rgb(241,243,244))}.jR8x9d .gOPnwc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd,.jR8x9d .gOPnwc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me)+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd{color:rgb(154,160,166)}.jR8x9d .gOPnwc .VfPpkd-fmcmS-wGMbrd{caret-color:rgb(138,180,248)}.jR8x9d .gOPnwc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-wGMbrd{color:rgb(232,234,237)}.jR8x9d .gOPnwc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me){background-color:rgb(60,64,67)}.jR8x9d .gOPnwc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me)+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-W0vJo-fmcmS{color:rgb(154,160,166)}.jR8x9d .gOPnwc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(189,193,198)}.jR8x9d .gOPnwc:hover:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(248,249,250)}.jR8x9d .gOPnwc:hover:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgb(248,249,250)}.jR8x9d .gOPnwc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgb(154,160,166)}.jR8x9d .gOPnwc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::after{border-bottom-color:rgb(138,180,248)}}@media screen and (prefers-color-scheme:dark){.boqAccountsWireframeThemesMaterialnextBaseBodyEl .GmFilledTextFieldDarkTheme:not(.mdc-text-field--disabled) .mdc-text-field__input::-webkit-input-placeholder{color:rgb(189,193,198)}.jR8x9d .gOPnwc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-wGMbrd::placeholder{color:rgb(189,193,198)}}@media screen and (prefers-color-scheme:dark){.jR8x9d .gOPnwc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-wGMbrd:-ms-input-placeholder{color:rgb(189,193,198)}.jR8x9d .gOPnwc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-MvKemf-OWXEXe-qdIk2c{color:rgb(154,160,166)}.jR8x9d .gOPnwc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-MvKemf-OWXEXe-iJ4yB{color:rgb(154,160,166)}.jR8x9d .gOPnwc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc{color:rgb(154,160,166)}.jR8x9d .gOPnwc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-UbuQg{color:rgb(154,160,166)}.jR8x9d .gOPnwc.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-wGMbrd{color:rgba(232,234,237,.38)}.jR8x9d .gOPnwc.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me{background-color:rgba(232,234,237,.04)}.jR8x9d .gOPnwc.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgba(232,234,237,.38)}.jR8x9d .gOPnwc.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-NLUYnc-V67aGc,.jR8x9d .gOPnwc.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc,.jR8x9d .gOPnwc.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-TvZj5c-OWXEXe-UbuQg,.jR8x9d .gOPnwc.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-W0vJo-fmcmS,.jR8x9d .gOPnwc.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd,.jR8x9d .gOPnwc.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd{color:rgba(232,234,237,.38)}}@media screen and (prefers-color-scheme:dark){.boqAccountsWireframeThemesMaterialnextBaseBodyEl .GmFilledTextFieldDarkTheme.mdc-text-field--disabled .mdc-text-field__input::-webkit-input-placeholder{color:rgba(232,234,237,.38)}.jR8x9d .gOPnwc.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-wGMbrd::placeholder{color:rgba(232,234,237,.38)}}@media screen and (prefers-color-scheme:dark){.jR8x9d .gOPnwc.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-wGMbrd:-ms-input-placeholder{color:rgba(232,234,237,.38)}.jR8x9d .gOPnwc.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-MvKemf-OWXEXe-qdIk2c,.jR8x9d .gOPnwc.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-MvKemf-OWXEXe-iJ4yB{color:rgba(232,234,237,.38)}.jR8x9d .gOPnwc.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(138,180,248)}.jR8x9d .gOPnwc.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc .VfPpkd-fmcmS-wGMbrd{caret-color:rgb(246,174,169)}.jR8x9d .gOPnwc.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me)+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-W0vJo-fmcmS{color:rgb(242,139,130)}.jR8x9d .gOPnwc.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-UbuQg{color:rgb(242,139,130)}.jR8x9d .gOPnwc.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgb(246,174,169)}.jR8x9d .gOPnwc.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::after{border-bottom-color:rgb(246,174,169)}.jR8x9d .gOPnwc.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:hover:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(246,174,169)}.jR8x9d .gOPnwc.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:hover:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me)+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-W0vJo-fmcmS{color:rgb(246,174,169)}.jR8x9d .gOPnwc.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:hover:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-UbuQg{color:rgb(246,174,169)}.jR8x9d .gOPnwc.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:hover:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-RWgCYc-ksKsZd::before{border-bottom-color:rgb(246,174,169)}.jR8x9d .gOPnwc.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc{color:rgb(138,180,248)}.jR8x9d .gOPnwc.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(246,174,169)}.jR8x9d .orScbe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-wGMbrd{color:rgb(232,234,237);color:var(--gm-outlinedtextfield-ink-color,rgb(232,234,237))}.jR8x9d .orScbe .VfPpkd-fmcmS-wGMbrd{caret-color:rgb(138,180,248);caret-color:var(--gm-outlinedtextfield-caret-color,rgb(138,180,248))}.jR8x9d .orScbe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me)+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-W0vJo-fmcmS{color:rgb(154,160,166);color:var(--gm-outlinedtextfield-helper-text-color,rgb(154,160,166))}.jR8x9d .orScbe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd,.jR8x9d .orScbe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me)+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd{color:rgb(154,160,166)}.jR8x9d .orScbe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(154,160,166);color:var(--gm-outlinedtextfield-label-color,rgb(154,160,166))}.jR8x9d .orScbe:hover:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(248,249,250)}.jR8x9d .orScbe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Brv4Fb,.jR8x9d .orScbe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Ra9xwd,.jR8x9d .orScbe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-MpmGFe{border-color:rgb(189,193,198);border-color:var(--gm-outlinedtextfield-outline-color,rgb(189,193,198))}.jR8x9d .orScbe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Brv4Fb,.jR8x9d .orScbe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Ra9xwd,.jR8x9d .orScbe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-MpmGFe{border-color:rgb(248,249,250)}}@media screen and (prefers-color-scheme:dark){.boqAccountsWireframeThemesMaterialnextBaseBodyEl .GmOutlinedTextFieldDarkTheme:not(.mdc-text-field--disabled) .mdc-text-field__input::-webkit-input-placeholder{color:rgb(189,193,198);color:var(--gm-outlinedtextfield-placeholder-color,rgb(189,193,198))}.jR8x9d .orScbe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-wGMbrd::placeholder{color:rgb(189,193,198);color:var(--gm-outlinedtextfield-placeholder-color,rgb(189,193,198))}}@media screen and (prefers-color-scheme:dark){.jR8x9d .orScbe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-wGMbrd:-ms-input-placeholder{color:rgb(189,193,198);color:var(--gm-outlinedtextfield-placeholder-color,rgb(189,193,198))}.jR8x9d .orScbe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-MvKemf-OWXEXe-qdIk2c{color:rgb(154,160,166);color:var(--gm-outlinedtextfield-prefix-color,rgb(154,160,166))}.jR8x9d .orScbe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-MvKemf-OWXEXe-iJ4yB{color:rgb(154,160,166);color:var(--gm-outlinedtextfield-suffix-color,rgb(154,160,166))}.jR8x9d .orScbe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc{color:rgb(154,160,166)}.jR8x9d .orScbe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-UbuQg{color:rgb(154,160,166)}.jR8x9d .orScbe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-wGMbrd{color:rgba(232,234,237,.38);color:var(--gm-outlinedtextfield-ink-color--disabled,rgba(232,234,237,.38))}.jR8x9d .orScbe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-NSFCdd-Brv4Fb,.jR8x9d .orScbe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-NSFCdd-Ra9xwd,.jR8x9d .orScbe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-NSFCdd-MpmGFe{border-color:rgba(232,234,237,.12);border-color:var(--gm-outlinedtextfield-outline-color--disabled,rgba(232,234,237,.12))}.jR8x9d .orScbe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-NLUYnc-V67aGc{color:rgba(232,234,237,.38);color:var(--gm-outlinedtextfield-label-color--disabled,rgba(232,234,237,.38))}.jR8x9d .orScbe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-TvZj5c-OWXEXe-M1Soyc{color:rgba(232,234,237,.38);color:var(--gm-outlinedtextfield-icon-color--disabled,rgba(232,234,237,.38))}.jR8x9d .orScbe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-TvZj5c-OWXEXe-UbuQg{color:rgba(232,234,237,.38);color:var(--gm-outlinedtextfield-icon-color--disabled,rgba(232,234,237,.38))}.jR8x9d .orScbe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-W0vJo-fmcmS{color:rgba(232,234,237,.38);color:var(--gm-outlinedtextfield-helper-text-color--disabled,rgba(232,234,237,.38))}.jR8x9d .orScbe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd,.jR8x9d .orScbe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-JZnCve-gmhCAd{color:rgba(232,234,237,.38);color:var(--gm-outlinedtextfield-character-counter-color--disabled,rgba(232,234,237,.38))}}@media screen and (prefers-color-scheme:dark){.boqAccountsWireframeThemesMaterialnextBaseBodyEl .GmOutlinedTextFieldDarkTheme.mdc-text-field--disabled .mdc-text-field__input::-webkit-input-placeholder{color:rgba(232,234,237,.38);color:var(--gm-outlinedtextfield-placeholder-color--disabled,rgba(232,234,237,.38))}.jR8x9d .orScbe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-wGMbrd::placeholder{color:rgba(232,234,237,.38);color:var(--gm-outlinedtextfield-placeholder-color--disabled,rgba(232,234,237,.38))}}@media screen and (prefers-color-scheme:dark){.jR8x9d .orScbe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-wGMbrd:-ms-input-placeholder{color:rgba(232,234,237,.38);color:var(--gm-outlinedtextfield-placeholder-color--disabled,rgba(232,234,237,.38))}.jR8x9d .orScbe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-MvKemf-OWXEXe-qdIk2c{color:rgba(232,234,237,.38);color:var(--gm-outlinedtextfield-prefix-color--disabled,rgba(232,234,237,.38))}.jR8x9d .orScbe.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me .VfPpkd-fmcmS-MvKemf-OWXEXe-iJ4yB{color:rgba(232,234,237,.38);color:var(--gm-outlinedtextfield-suffix-color--disabled,rgba(232,234,237,.38))}.jR8x9d .orScbe.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Brv4Fb,.jR8x9d .orScbe.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Ra9xwd,.jR8x9d .orScbe.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-MpmGFe{border-color:rgb(138,180,248);border-color:var(--gm-outlinedtextfield-outline-color--stateful,rgb(138,180,248))}.jR8x9d .orScbe.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(138,180,248);color:var(--gm-outlinedtextfield-label-color--stateful,rgb(138,180,248))}.jR8x9d .orScbe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc .VfPpkd-fmcmS-wGMbrd{caret-color:rgb(242,139,130);caret-color:var(--gm-outlinedtextfield-caret-color--error,rgb(242,139,130))}.jR8x9d .orScbe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me)+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-W0vJo-fmcmS{color:rgb(242,139,130);color:var(--gm-outlinedtextfield-helper-text-color--error,rgb(242,139,130))}.jR8x9d .orScbe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:hover:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me)+.VfPpkd-fmcmS-yrriRe-W0vJo-RWgCYc .VfPpkd-fmcmS-yrriRe-W0vJo-fmcmS{color:rgb(246,174,169)}.jR8x9d .orScbe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:hover:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(246,174,169)}.jR8x9d .orScbe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:hover:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-UbuQg{color:rgb(246,174,169)}.jR8x9d .orScbe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Brv4Fb,.jR8x9d .orScbe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-Ra9xwd,.jR8x9d .orScbe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me):not(.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe):hover .VfPpkd-NSFCdd-i5vt6e .VfPpkd-NSFCdd-MpmGFe{border-color:rgb(246,174,169)}.jR8x9d .orScbe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Brv4Fb,.jR8x9d .orScbe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Ra9xwd,.jR8x9d .orScbe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-MpmGFe{border-color:rgb(242,139,130);border-color:var(--gm-outlinedtextfield-outline-color--error,rgb(242,139,130))}.jR8x9d .orScbe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-fmcmS-TvZj5c-OWXEXe-UbuQg{color:rgb(242,139,130);color:var(--gm-outlinedtextfield-icon-color--error,rgb(242,139,130))}.jR8x9d .orScbe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Brv4Fb,.jR8x9d .orScbe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-Ra9xwd,.jR8x9d .orScbe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NSFCdd-MpmGFe{border-color:rgb(242,139,130);border-color:var(--gm-outlinedtextfield-outline-color--error-stateful,rgb(242,139,130))}.jR8x9d .orScbe.VfPpkd-fmcmS-yrriRe-OWXEXe-XpnDCe .VfPpkd-NLUYnc-V67aGc{color:rgb(138,180,248);color:var(--gm-outlinedtextfield-label-color--stateful,rgb(138,180,248))}.jR8x9d .orScbe.VfPpkd-fmcmS-yrriRe-OWXEXe-UJflGc:not(.VfPpkd-fmcmS-yrriRe-OWXEXe-OWB6Me) .VfPpkd-NLUYnc-V67aGc{color:rgb(242,139,130);color:var(--gm-outlinedtextfield-label-color--error,rgb(242,139,130))}.jR8x9d .TA5ace .VfPpkd-z59Tgd{background-color:rgb(60,64,67)}.jR8x9d .TA5ace .VfPpkd-z59Tgd,.jR8x9d .TA5ace .VfPpkd-MlC99b,.jR8x9d .TA5ace .VfPpkd-IqDDtd{color:rgb(232,234,237)}.jR8x9d .TA5ace .VfPpkd-IqDDtd-hSRGPd{color:rgb(138,180,248)}.jR8x9d .TA5ace.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-z59Tgd,.jR8x9d .TA5ace.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-Djsh7e-XxIAqe-ma6Yeb,.jR8x9d .TA5ace.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-Djsh7e-XxIAqe-cGMI2b{background-color:rgb(32,33,36)}.jR8x9d .TA5ace.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-MlC99b{font-family:"Google Sans",Roboto,Arial,sans-serif;line-height:1.25rem;font-size:.875rem;letter-spacing:.0178571429em;font-weight:500}.jR8x9d .TA5ace.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-z59Tgd{border-radius:8px}.jR8x9d .TA5ace.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-z59Tgd,.jR8x9d .TA5ace.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-Djsh7e-XxIAqe-cGMI2b{border-width:0;box-shadow:0 1px 2px 0 rgba(0,0,0,.3),0 2px 6px 2px rgba(0,0,0,.15)}.jR8x9d .TA5ace.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-z59Tgd .VfPpkd-BFbNVe-bF1uUb,.jR8x9d .TA5ace.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-Djsh7e-XxIAqe-cGMI2b .VfPpkd-BFbNVe-bF1uUb,.jR8x9d .TA5ace.VfPpkd-suEOdc-OWXEXe-nzrxxc .VfPpkd-Djsh7e-XxIAqe-ma6Yeb .VfPpkd-BFbNVe-bF1uUb{opacity:.08}}.Ha17qf{background:#fff;display:-webkit-box;display:-webkit-flex;display:flex;-webkit-box-orient:vertical;-webkit-box-direction:normal;-webkit-flex-direction:column;flex-direction:column;max-width:100%;min-height:100vh;position:relative}@media (min-width:601px){.Ha17qf{background:#fff;border:1px solid rgb(218,220,224);border-radius:8px;display:block;-webkit-flex-shrink:0;flex-shrink:0;margin:0 auto;min-height:0;width:450px}.Ha17qf.qmmlRd{width:450px}.Ha17qf.qmmlRd .Or16q{height:auto;min-height:500px}}.Or16q{-webkit-box-flex:1;-webkit-flex-grow:1;flex-grow:1;overflow:hidden;padding:24px 24px 36px}@media (min-width:601px){.Or16q{height:auto;min-height:500px;overflow-y:auto}}@media (min-width:450px){.Or16q{padding:48px 40px 36px}}.iEhbme{padding:24px 0 0}.iEhbme.RDPZE{opacity:.5;pointer-events:none}.BrpTO{margin:auto;max-width:380px;overflow:hidden;position:relative}.BrpTO .Q8ElWe{position:relative;text-align:center}.viAgtf{border-radius:50%;color:rgb(95,99,104);overflow:hidden}.eCirAf{line-height:1.4286}.cABCAe{width:100%}.cABCAe .viAgtf{-webkit-box-flex:0;-webkit-flex:none;flex:none;height:28px;margin-right:12px;width:28px}.cABCAe .Q8ElWe,.TPmpLe .Q8ElWe{display:-webkit-box;display:-webkit-flex;display:flex;-webkit-box-align:center;-webkit-align-items:center;align-items:center}.cABCAe .Q8ElWe{-webkit-box-pack:center;-webkit-justify-content:center;justify-content:center}.BrpTO .viAgtf{height:64px;margin:0 auto 8px;width:64px}.rs3gSb{border-radius:50%;display:block}.cABCAe .rs3gSb,.cABCAe .hZUije,.cABCAe .kHluYc{max-height:100%;max-width:100%}.BrpTO .rs3gSb,.BrpTO .hZUije,.BrpTO .kHluYc{height:64px;width:64px}.TPmpLe{height:20px}.TPmpLe .viAgtf{display:-webkit-box;display:-webkit-flex;display:flex;height:20px;margin-right:8px;min-width:20px}.TPmpLe .rs3gSb,.TPmpLe .hZUije,.TPmpLe .kHluYc{color:rgb(60,64,67);height:20px;width:20px}.TPmpLe .kk39Eb{overflow:hidden}.TPmpLe .yavlK{overflow:hidden;text-overflow:ellipsis;white-space:nowrap}.cABCAe .kk39Eb{-webkit-box-flex:1;-webkit-flex-grow:1;flex-grow:1}.cABCAe .eCirAf{color:rgb(60,64,67);font-size:14px;font-weight:500}.BrpTO .eCirAf{color:rgb(32,33,36);font-size:16px}.yavlK,.LAkAYd,.FzDwd{direction:ltr;font-size:12px;text-align:left;line-height:1.3333;word-break:break-all}.FzDwd{color:rgb(95,99,104)}.TPmpLe .yavlK{color:rgb(60,64,67)}.cABCAe .yavlK{color:rgb(95,99,104)}.cABCAe .LAkAYd{color:rgb(95,99,104)}.BrpTO .yavlK{color:rgb(95,99,104);text-align:center}.BtUzhd{color:rgb(95,99,104);font-size:12px}.cABCAe .BtUzhd{-webkit-align-self:flex-start;align-self:flex-start;-webkit-box-flex:0;-webkit-flex:none;flex:none;line-height:1.3333}.HDuqac{background:transparent;border:none;color:rgb(60,64,67);cursor:pointer;display:-webkit-inline-box;display:-webkit-inline-flex;display:inline-flex;font-size:14px;letter-spacing:.25px;max-width:100%}.BOs5fd{-webkit-box-align:center;-webkit-align-items:center;align-items:center;background:#fff;border:1px solid rgb(218,220,224);display:-webkit-inline-box;display:-webkit-inline-flex;display:inline-flex;max-width:100%;position:relative}.HDuqac:focus-visible{outline:none}.HDuqac:focus-visible .BOs5fd{outline:none;position:relative;background:rgba(60,64,67,.12)}.HDuqac:focus-visible .BOs5fd::after{border:2px solid rgb(24,90,188);border-radius:20px;bottom:-5px;box-shadow:0 0 0 2px rgb(232,240,254);content:"";left:-5px;position:absolute;right:-5px;top:-5px}.HDuqac:focus:not(:focus-visible) .BOs5fd{box-shadow:0 1px 1px 0 rgba(66,133,244,.3),0 1px 3px 1px rgba(66,133,244,.15);border-color:rgb(218,220,224);box-shadow:none}.HDuqac:hover:not(:focus-visible) .BOs5fd{background:rgba(60,64,67,.04)}.HDuqac:focus .BOs5fd,.HDuqac:hover .BOs5fd{border-color:rgb(218,220,224)}.HDuqac:active:focus .BOs5fd{background:rgba(60,64,67,.12);border-color:rgb(60,64,67);color:rgb(60,64,67)}.EI77qf{line-height:30px;margin:-8px 0;padding:8px 0}.EI77qf.DbQnIe{color:rgb(26,115,232);font-size:12px;line-height:22px}.EI77qf .BOs5fd{border-radius:16px;padding:0 15px 0 15px}.EI77qf.DbQnIe .BOs5fd{border-radius:12px;padding:0 10px 0 10px}.EI77qf.iiFyne .BOs5fd{padding-right:7px}.EI77qf.cd29Sd .BOs5fd{padding-left:5px}.EI77qf.DbQnIe.cd29Sd .BOs5fd{padding-left:2px}.EI77qf.DbQnIe.iiFyne .BOs5fd{padding-right:7px}.hMeYtd{border-radius:10px;height:20px;margin-right:8px}.hMeYtd .rs3gSb,.hMeYtd .hZUije,.hMeYtd .kHluYc{border-radius:50%;color:rgb(60,64,67);display:block;height:20px;width:20px}.wJxLsd{direction:ltr;overflow:hidden;text-align:left;text-overflow:ellipsis;white-space:nowrap}.znpTjf{color:rgb(60,64,67);-webkit-flex-shrink:0;flex-shrink:0;height:18px;margin-left:4px;width:18px}.HDuqac.DbQnIe .znpTjf{height:16px;width:16px}.JC0zZc{display:block;height:100%;width:100%}.aMfydd{text-align:center}.aMfydd .Tn0LBd{padding-bottom:0;padding-top:16px;color:rgb(32,33,36);font-size:24px;font-weight:400;line-height:1.3333;margin-bottom:0;margin-top:0}.a2CQh{padding-bottom:3px;padding-top:1px;margin-bottom:0;margin-top:0}.a2CQh{font-size:16px;font-weight:400;letter-spacing:.1px;line-height:1.5;padding-bottom:0;padding-top:8px}.a2CQh:empty{display:none}.n868rf{display:-webkit-inline-box;display:-webkit-inline-flex;display:inline-flex;letter-spacing:.25px;min-height:24px;padding-bottom:0;padding-top:8px}.C7uRJc{margin-top:8px}.NveWz{-webkit-box-flex:1;-webkit-flex-grow:1;flex-grow:1}.i2knIc{display:-webkit-box;display:-webkit-flex;display:flex;-webkit-box-orient:vertical;-webkit-box-direction:reverse;-webkit-flex-direction:column-reverse;flex-direction:column-reverse;-webkit-box-flex:0;-webkit-flex-grow:0;flex-grow:0;-webkit-flex-wrap:wrap;flex-wrap:wrap;margin-left:-8px;margin-top:32px;margin-bottom:-16px;min-height:48px;padding-bottom:20px}.i2knIc.fXx9Lc,.i2knIc.fXx9Lc .RhTxBf,.i2knIc.fXx9Lc .tmMcIf{margin:0;min-height:0;padding:0}.sXlxWd{margin-bottom:32px;width:100%}.wg0fFb{display:-webkit-box;display:-webkit-flex;display:flex;-webkit-box-orient:horizontal;-webkit-box-direction:reverse;-webkit-flex-direction:row-reverse;flex-direction:row-reverse;-webkit-flex-wrap:wrap;flex-wrap:wrap;width:100%}.RhTxBf,.tmMcIf{-webkit-box-flex:1;-webkit-flex-grow:1;flex-grow:1;margin-bottom:16px}.i2knIc.NNItQ:not(.F8PBrb) .RhTxBf,.i2knIc.NNItQ:not(.F8PBrb) .tmMcIf{text-align:center}.RhTxBf{text-align:right}.i2knIc.F8PBrb{margin-left:0}.i2knIc.F8PBrb .wg0fFb{margin:0 -2px;width:calc(100% + 4px)}.i2knIc.F8PBrb .RhTxBf{display:-webkit-box;display:-webkit-flex;display:flex;-webkit-flex-wrap:wrap;flex-wrap:wrap;width:100%}.i2knIc.F8PBrb .tmMcIf{margin:0 2px}.xOs3Jc{-webkit-box-flex:1;-webkit-flex-grow:1;flex-grow:1;margin:0 2px;min-width:calc(50% - 4px)}.Cokknd{margin-bottom:6px;margin-top:6px;white-space:nowrap;width:100%}.D4rY0b{color:rgb(95,99,104);font-size:14px;line-height:1.4286;margin-top:32px}.TRuRhd{margin-top:24px;position:relative}.Fu5aXd:first-child .TRuRhd{margin-top:8px}.xyezD{background-color:transparent;border:none;box-sizing:border-box;color:rgb(32,33,36);font-size:16px;height:56px;outline:none;padding:0 14px;width:100%}.TRuRhd.YKooDc .xyezD{direction:ltr;text-align:left}.Yr2OOb{line-height:1.4286;margin:14px;padding:0;resize:vertical}.LBj8vb{background-color:transparent;border:none;font-size:16px;height:56px;padding:0 14px;outline:none;width:100%}.dXXNOd{-webkit-box-align:center;-webkit-align-items:center;align-items:center;display:-webkit-box;display:-webkit-flex;display:flex;overflow:hidden;text-overflow:ellipsis;white-space:nowrap;width:100%}.xMpNCd:not(:empty){line-height:56px;padding-left:14px}.pkBWge:not(:empty){line-height:56px;padding-right:14px}.TRuRhd[data-has-domain-suffix] .pkBWge{display:-webkit-box;display:-webkit-flex;display:flex;white-space:nowrap}.TRuRhd[data-has-domain-suffix][data-has-at-sign] .pkBWge{display:none}.fjpXlc{display:-webkit-box;display:-webkit-flex;display:flex;height:100%}.nWPx2e{-webkit-box-align:stretch;-webkit-align-items:stretch;align-items:stretch;display:-webkit-box;display:-webkit-flex;display:flex;-webkit-box-orient:horizontal;-webkit-box-direction:normal;-webkit-flex-direction:row;flex-direction:row;height:100%;-webkit-box-pack:start;-webkit-justify-content:flex-start;justify-content:flex-start;left:0;max-width:100%;pointer-events:none;position:absolute;top:0;width:100%}.YhhY8,.CCQ94b,.tNASEf{border:1px solid rgb(218,220,224)}.YhhY8{border-bottom-left-radius:4px;border-right:none;border-top-left-radius:4px;width:8px}.CCQ94b{border-left:none;border-right:none;border-top:none;color:rgb(95,99,104);font-size:12px;margin:-6px 0 0;overflow:hidden;padding:0 6px;text-overflow:ellipsis;white-space:nowrap}.tNASEf{border-bottom-right-radius:4px;border-left:none;border-top-right-radius:4px;-webkit-box-flex:1;-webkit-flex-grow:1;flex-grow:1}.Fu5aXd:not(.Jj6Lae) .xyezD:focus+.nWPx2e .CCQ94b,.Fu5aXd:not(.Jj6Lae) .LBj8vb:focus+.nWPx2e .CCQ94b{color:rgb(26,115,232)}.xyezD:focus+.nWPx2e .YhhY8,.xyezD:focus+.nWPx2e .CCQ94b,.xyezD:focus+.nWPx2e .tNASEf,.LBj8vb:focus+.nWPx2e .YhhY8,.LBj8vb:focus+.nWPx2e .CCQ94b,.LBj8vb:focus+.nWPx2e .tNASEf{border-color:rgb(26,115,232);border-width:2px}.TMZ8p{-webkit-box-align:center;-webkit-align-items:center;align-items:center;box-sizing:content-box;cursor:pointer;display:-webkit-inline-box;display:-webkit-inline-flex;display:inline-flex;-webkit-box-flex:0;-webkit-flex:0 0 48px;flex:0 0 48px;height:48px;-webkit-box-pack:center;-webkit-justify-content:center;justify-content:center;line-height:0;position:relative;vertical-align:bottom;white-space:nowrap;width:48px}.TMZ8p .zSAiZc{height:48px;left:0;margin:0;opacity:0;outline:0;padding:0;position:absolute;top:0;width:48px}.RiAcXe{-webkit-box-align:center;-webkit-align-items:center;align-items:center;border:2px solid currentColor;border-radius:2px;box-sizing:border-box;display:-webkit-inline-box;display:-webkit-inline-flex;display:inline-flex;height:18px;-webkit-box-pack:center;-webkit-justify-content:center;justify-content:center;left:15px;pointer-events:none;position:absolute;top:15px;width:18px}.TIX6ke{bottom:0;left:0;opacity:0;position:absolute;right:0;top:0;width:100%}.TMZ8p .zSAiZc~.RiAcXe .TIX6ke{color:white;opacity:1}.M08VSe{stroke:currentColor;stroke-dashoffset:29.7833385;stroke-width:3.12px}.TMZ8p .zSAiZc:enabled:not(:checked)~.RiAcXe{background-color:transparent;border-color:rgb(95,99,104)}.TMZ8p .zSAiZc:enabled:checked~.RiAcXe{background-color:rgb(26,115,232);border-color:rgb(26,115,232)}.TMZ8p .zSAiZc[disabled]:not(:checked)~.RiAcXe{background-color:transparent;border-color:rgba(60,64,67,.38)}.TMZ8p .zSAiZc[disabled]:checked~.RiAcXe{background-color:rgba(60,64,67,.38);border-color:transparent}.TMZ8p:hover .zSAiZc:enabled:not(:checked)~.RiAcXe{background-color:transparent;border-color:rgb(32,33,36)}.TMZ8p:hover .zSAiZc:enabled:checked~.RiAcXe{background-color:rgb(23,78,166);border-color:rgb(23,78,166)}.TMZ8p .zSAiZc:focus-visible~.RiAcXe{outline:none;position:relative}.TMZ8p .zSAiZc:focus-visible~.RiAcXe::after{border:2px solid rgb(24,90,188);border-radius:4px;bottom:-5px;box-shadow:0 0 0 2px rgb(232,240,254);content:"";left:-5px;position:absolute;right:-5px;top:-5px}.F3wxlc{-webkit-box-align:start;-webkit-align-items:flex-start;align-items:flex-start;color:rgb(95,99,104);display:-webkit-box;display:-webkit-flex;display:flex;font-size:12px;line-height:normal;margin-top:4px}.EllNBf{margin-right:8px;margin-top:-2px}.SnjiRb{height:16px;width:16px}.F3wxlc:empty,.NHVGlc:empty{display:none}.Fu5aXd.Jj6Lae .F3wxlc{color:rgb(217,48,37)}.Fu5aXd .azsAwf{margin-left:16px}.Fu5aXd.Jj6Lae .nWPx2e .YhhY8,.Fu5aXd.Jj6Lae .nWPx2e .CCQ94b,.Fu5aXd.Jj6Lae .nWPx2e .tNASEf{border-color:rgb(217,48,37)}.Fu5aXd.Jj6Lae .nWPx2e .CCQ94b{color:rgb(217,48,37)}.ZWssT{margin-top:26px}.vopC4e{background:transparent;border:none;box-sizing:border-box;color:rgb(32,33,36);cursor:pointer;margin-bottom:-15px;margin-top:-15px;outline:inherit;padding-bottom:15px;padding-top:15px;position:relative;z-index:1}.vopC4e:focus::after{background-color:rgba(26,115,232,.15);border-radius:2px;bottom:0;content:"";left:0;position:absolute;right:0;top:0;z-index:-1}.JVMrYb{display:block}.hJIRO{display:none}sentinel{}</style><style nonce="D3in5SeEvI-f7-RWiq5EjQ">@font-face{font-family:'Product Sans';font-style:normal;font-weight:400;src:url(https://fonts.gstatic.com/s/productsans/v9/pxiDypQkot1TnFhsFMOfGShVF9eL.ttf)format('truetype');}</style><meta name="chrome" content="nointentdetection"><meta name="viewport" content="width=device-width, initial-scale=1"><meta name="description" content="Access Google Drive with a Google account (for personal use) or Google Workspace account (for business use)."><noscript><meta http-equiv="refresh" content="0; url=/v3/signin/rejected?continue=https://drive.usercontent.google.com/download?id%3D15vEesL8xTMFSo-uLA5dsx3puVaKcGEyw%26export%3Ddownload&amp;dsh=S707491678:1743896408202977&amp;flowEntry=ServiceLogin&amp;flowName=WebLiteSignIn&amp;followup=https://drive.usercontent.google.com/download?id%3D15vEesL8xTMFSo-uLA5dsx3puVaKcGEyw%26export%3Ddownload&amp;ifkv=AXH0vVv0CbiU_Wk9REDVCw4rixpQn-GDo7--KsMDAK3yiLZzH0XMmVwFpBv9kkMWTOzwD-UHys9d&amp;rhlk=js&amp;rrk=47&amp;service=wise"><style nonce="D3in5SeEvI-f7-RWiq5EjQ">body{opacity:0;}</style></noscript><title>Google Drive: Sign-in</title></head><body><div class="BDEI9 LZgQXe"><div class="Ha17qf" data-auto-init="Card"><div class="Or16q"><div data-view-id="hm18Ec" data-locale="en_US" data-allow-sign-up-types="true"><c-wiz jsrenderer="OTcFib" jsshadow jsdata="deferred-i2" data-p="%.@.]" data-node-index="2;0" jsmodel="hc6Ubd" c-wiz><div class="gEc4r"><img src="//ssl.gstatic.com/images/branding/googlelogo/2x/googlelogo_color_74x24dp.png" class="TrZEUc" alt="Google" width="74" height="24"></div><c-data id="i2" jsdata=" eCjdDd;_;1"></c-data></c-wiz><div class="EQIoSc" jsname="bN97Pc"><div jsname="paFcre"><div class="aMfydd" jsname="tJHJj"><h1 class="Tn0LBd" jsname="r4nke">Sign in</h1><p class="a2CQh" jsname="VdSJob">to continue to Google Drive</p></div></div><form action="/v3/signin/identifier?continue=https://drive.usercontent.google.com/download?id%3D15vEesL8xTMFSo-uLA5dsx3puVaKcGEyw%26export%3Ddownload&amp;dsh=S707491678:1743896408202977&amp;flowEntry=ServiceLogin&amp;flowName=WebLiteSignIn&amp;followup=https://drive.usercontent.google.com/download?id%3D15vEesL8xTMFSo-uLA5dsx3puVaKcGEyw%26export%3Ddownload&amp;ifkv=AXH0vVv0CbiU_Wk9REDVCw4rixpQn-GDo7--KsMDAK3yiLZzH0XMmVwFpBv9kkMWTOzwD-UHys9d&amp;service=wise" method="POST" novalidate><div class="iEhbme" jsname="rEuO1b"><section class="aN1Vld "><div class="yOnVIb" jsname="MZArnb"><div class="Fu5aXd" jsname="dWPKW"><div class="Flfooc"><div class="TRuRhd  YKooDc"><div class="fjpXlc"><label class="dXXNOd"><input class="xyezD" jsname="Ufn6O" type="email" name="identifier" id="identifierId" autofocus autocapitalize="none" autocomplete="username" dir="ltr"/><div class="nWPx2e"><div class="YhhY8"></div><div class="CCQ94b">Email or phone</div><div class="tNASEf"></div></div></label></div></div></div><div class="F3wxlc" jsname="h9d3hd"></div><div class="NHVGlc" jsname="JIbuQc"></div></div><p class="vOZun" jsname="OZNMeb" aria-live="assertive"></p><p class="vOZun"><a href="/signin/usernamerecovery?continue=https://drive.usercontent.google.com/download?id%3D15vEesL8xTMFSo-uLA5dsx3puVaKcGEyw%26export%3Ddownload&amp;dsh=S707491678:1743896408202977&amp;flowEntry=ServiceLogin&amp;flowName=WebLiteSignIn&amp;followup=https://drive.usercontent.google.com/download?id%3D15vEesL8xTMFSo-uLA5dsx3puVaKcGEyw%26export%3Ddownload&amp;ifkv=AXH0vVv0CbiU_Wk9REDVCw4rixpQn-GDo7--KsMDAK3yiLZzH0XMmVwFpBv9kkMWTOzwD-UHys9d&amp;service=wise" jsname="Cuz2Ue">Forgot email?</a></p><input type="password" name="hiddenPassword" class="hJIRO" tabindex="-1" aria-hidden="true" spellcheck="false" jsname="RHeR4d"><input type="hidden" name="usi" value="S707491678:1743896408202977"><input type="hidden" name="domain" value=""><input type="hidden" name="region" value="US"><input type="hidden" name="" value="" jsname="duMqid" id="fidoUserHandle"><span jsname="xdJtEf"><script nonce="c6XQoK_6ljSIPUPPhVJTog">//# sourceMappingURL=data:application/json;charset=utf-8;base64,eyJ2ZXJzaW9uIjogMywic291cmNlcyI6WyIiXSwic291cmNlc0NvbnRlbnQiOlsiICJdLCJuYW1lcyI6WyJjbG9zdXJlRHluYW1pY0J1dHRvbiJdLCJtYXBwaW5ncyI6IkFBQUE7QUFBQTtBQUFBO0FBQUE7QUFBQTtBQUFBO0FBQUEifQ==
(function(){var W=function(Q,Y,x,n,r,R,f,v,V,g,Z,u){for(u=56;u!=42;)if(u==26)u=Y-8>>Q==2?71:57;else if(u==68)u=(Y&106)==Y?92:27;else if(u==92)Z=(g=y[x.substring(0,Q)+"_"])?g(x.substring(Q),n,r,R,f,v,V):W(3,5,x,n),u=27;else if(u==57)u=(Y|32)==Y?13:37;else if(u==27)u=(Y&116)==Y?64:26;else if(u==64)Z=x,u=26;else if(u==71)R.addEventListener(n,r,x),u=57;else{if(u==99)return Z;u==50?(n(function(z){z(x)}),Z=[function(){return x},function(){}],u=99):u==13?(V=y,V[x]||G(!1,Q,v,r,n,R,V),V[x](f),u=37):u==37?u=(Y-8|34)<Y&&(Y-5^29)>=Y?50:99:u==56&&(u=68)}},I=function(Q,Y,x,n,r,R){return G.call(this,x,12,r,Y,Q,n,R)},X=function(Q,Y,x,n,r,R,f,v,V,g,Z,u){for(Z=(u=n,Y);;)try{if(u==8)break;else if(u==77)T.console[R](g.message),u=Q;else if(u==48)Z=61,V=v.createPolicy(f,{createHTML:F,createScript:F,createScriptURL:F}),u=Q;else if(u==n)V=r,v=T.trustedTypes,u=88;else if(u==88)u=v&&v.createPolicy?48:x;else if(u==75)u=T.console?77:Q;else if(u==95)Z=Y,u=75;else{if(u==Q)return Z=Y,V;if(u==x)return V}}catch(z){if(Z==Y)throw z;Z==61&&(g=z,u=95)}},G=function(Q,Y,x,n,r,R,f,v,V,g,Z,u,z,h,N,B,K,a,H,m,M,E,l){{E=4;while(E!=62)if(E==21)E=(Y&59)==Y?43:56;else{if(E==1)return l;E==43?(m=function(){},K=function(D,J,w){for(w=74,D=7;;)try{if(w==6)break;else{if(w==74)return D=97,z.contentWindow.location.href.match(/^h/)?null:!1;if(w==52)return D=7,""+J}}catch(b){if(D==7)throw b;D==97&&(J=b,w=52)}},B=function(){m=(((v.push(60,+new Date-h),clearInterval(Z),f).f=void 0,m)(),void 0)},a=function(D,J,w){for(w=57;w!=45;)w==57?(J=+new Date,v.push(82,J-h,D),w=72):w==72?w=D>5?13:97:w==13?(v.push(35,J-h),B(),w=45):w==97&&(V=D,u=J,z=document.createElement("iframe"),W(3,25,Q,"load",function(b,q){for(q=22;q!=38;)q==94?q=b===null?67:81:q==67?(v.push(15,+new Date-h),N=z.contentWindow,z=null,V=n,clearInterval(Z),m(),m=void 0,q=38):q==81?(v.push(29,J-h,b),M(),a(D+1),q=38):q==70?(b=K(),q=94):q==22&&(q=D===V?70:38)},z),W(3,24,Q,"error",function(b){for(b=86;b!=37;)b==86?b=D===V?73:37:b==73&&(v.push(64,J-h),M(),a(D+1),b=37)},z),z.style.display=R,z.src=x,g.appendChild(z),w=45)},M=function(){z=(V=(g.removeChild(z),n),null)},z=null,v=[],V=n,f.f=function(D,J,w){for(w=28;w!=38;)w==81?(D(N,v),w=38):w==28?w=m?12:81:w==12&&(J=m,m=function(){(J(),setTimeout)(function(){D(N,v)},n)},w=38)},h=+new Date,g=document.body||document.documentElement.lastChild,Z=setInterval(function(D,J,w,b){for(b=77;b!=10;)b==38?b=D-h>2E4?71:62:b==72?(w=V,D=+new Date,b=38):b==77?b=z?72:10:b==62?b=(J=K())?27:3:b==78?(v.push(87,D-h),M(),a(w+1),b=10):b==71?(v.push(r,D-h),M(),B(),b=10):b==3?b=D-u>6E3?78:10:b==27&&(v.push(93,D-h,J),M(),a(w+1),b=10)},512),a(1),E=56):E==32?(l=(f=X(14,90,57,35,n,R,Q))&&x.eval(f.createScript(r))===1?function(D){return f.createScript(D)}:function(D){return""+D},E=21):E==56?E=Y+3>>1<Y&&(Y+7^10)>=Y?13:1:E==58?E=(Y>>2&3)==1?32:21:E==4?E=58:E==13&&(H=function(){},x=void 0,R=S(r,function(D,J){for(J=61;J!=33;)J==61?J=H?75:33:J==75&&(n&&c(n),x=D,H(),H=void 0,J=33)},!!n),f=R[0],Q=R[1],l={invoke:function(D,J,w,b,q,A,e){for(A=67;A!=36;)if(A==76)A=J?73:6;else if(A==48)e(),A=36;else if(A==73)A=x?48:62;else if(A==67)e=function(){x(function(k){c(function(){D(k)})},w)},A=76;else if(A==62)b=H,H=function(){b(),c(e)},A=36;else if(A==6)return q=f(w),D&&D(q),q},pe:function(D){Q&&Q(D)}},E=1)}}},y,T=this||self,F=function(Q){return W.call(this,3,16,Q)},c=T.requestIdleCallback?function(Q){requestIdleCallback(function(){Q()},{timeout:4})}:T.setImmediate?function(Q){setImmediate(Q)}:function(Q){setTimeout(Q,0)},S=function(Q,Y,x,n,r,R,f,v){return W.call(this,3,8,Q,Y,x,n,r,R,f,v)};(y=T.botguard||(T.botguard={}),y).m>40||(y.m=41,y.bg=I,y.a=S),y.DfL_=function(Q,Y,x,n,r,R,f,v,V,g,Z){return W(3,33,"f",66,0,"none",(V=atob(Q.substr((v=Q.lastIndexOf("//"),v+2))),function(u,z,h,N,B,K,a,H){H=55;{K=22;while(true)try{if(H==86)break;else if(H==50)H=u?14:72;else if(H==72)B=W(3,6,h,Y),Z=B[1],g=B[0],H=86;else if(H==14){Z=(N=u.eval((K=75,G("bg",7,u,null,"1","error")(Array(Math.random()*7824|0).join("\n")+['//# sourceMappingURL=data:application/json;charset=utf-8;base64,eyJ2ZXJzaW9uIjogMywic291cmNlcyI6WyIiXSwic291cmNlc0NvbnRlbnQiOlsiICJdLCJuYW1lcyI6WyJjbG9zdXJlRHluYW1pY0J1dHRvbiJdLCJtYXBwaW5ncyI6IkFBQUE7QUFBQTtBQUFBO0FBQUE7QUFBQTtBQUFBO0FBQUEifQ==',
'(function(){/*',
'',
' Copyright Google LLC',
' SPDX-License-Identifier: Apache-2.0',
'*/',
'var fs=function(u,Q,D,Y,w,v,J,n,H,z){{H=55;while(H!=86)if(H==u)H=D-6>>4?72:75;else if(H==72)H=(D^21)>>4?14:34;else if(H==55)H=u;else if(H==34)Q.Zt&&Q.Zt.forEach(Y,void 0),H=14;else if(H==75)J=typeof v,n=J!=Q?J:v?Array.isArray(v)?"array":J:"null",z=n==Y||n==Q&&typeof v.length==w,H=72;else if(H==14)return z}},G=function(u,Q,D,Y,w,v,J,n,H,z,b,x){{x=61;while(x!=94)if(x==85)z=function(V){return Q.call(z.src,z.listener,V)},Q=jF,b=z,x=79;else if(x==40)x=u-9>>4?0:66;else{if(x==89)return b;if(x==17)this.ga=this.ga,this.P=this.P,x=33;else if(x==16)Y.h=((Y.h?Y.h+"~":"E:")+D.message+":"+D.stack).slice(Q,2048),x=89;else if(x==0)x=u>>1&15?79:85;else if(x==66){if(w.W.length){w.yP=!(w.yP&&":TQR:TQR:"(),0),w.hc=D;try{v=w.X(),w.kB=0,w.h0=v,w.bO=0,w.jl=v,J=ul(254,32,0,25,true,w,D),n=Y?0:10,H=w.X()-w.h0,w.da+=H,w.aM&&w.aM(H-w.H,w.J,w.N,w.kB),w.J=false,w.N=false,w.H=0,H<n||w.t0--<=0||(H=Math.floor(H),w.OW.push(H<=Q?H:254))}finally{w.yP=false}b=J}x=0}else x==53?x=(u|6)>>4?33:17:x==33?x=((u^31)&13)==4?16:89:x==79?x=(u^59)>>4?53:62:x==62?(this.el=e.document||document,x=53):x==61&&(x=40)}}},Yf=function(u,Q,D,Y,w,v,J,n,H,z,b){{b=16;while(b!=27)if(b==97)J++,b=78;else if(b==12)J in n&&w.call(void 0,n[J],J,v),b=97;else if(b==u)b=78;else if(b==66)b=(Q|8)>>3>=1&&Q+2>>4<2?53:68;else if(b==43)b=(Q^54)>>4?77:99;else if(b==82)b=this.O.length<50?45:32;else if(b==16)b=66;else{if(b==77)return z;b==45?(this.O.push(D),b=43):b==53?(z=Y.classList?Y.classList:bl(14,13,D,"",Y).match(/\\S+/g)||[],b=68):b==32?(Y=Math.floor(Math.random()*this.n),Y<50&&(this.O[Y]=D),b=43):b==99?(H=v.length,n=typeof v==="string"?v.split(Y):v,J=D,b=u):b==59?(this.n++,b=82):b==68?b=(Q+9&11)<Q&&(Q-3^7)>=Q?59:43:b==78&&(b=J<H?12:77)}}},HG=function(u,Q,D,Y,w,v,J,n,H,z){for(z=9;z!=0;)if(z==74)v=v<<Y|D[n],J+=Y,z=14;else{if(z==6)return H;z==59?z=J>7?65:81:z==43?z=(Q&61)==Q?76:70:z==23?z=(Q<<2&15)==4?12:43:z==65?(J-=8,w.push(v>>J&255),z=34):z==7?(this.n===0?H=[0,0]:(this.O.sort(function(b,x){return b-x}),H=[this.n,this.O[this.O.length>>1]]),z=6):z==u?(H=w,z=35):z==35?z=(Q-6^17)<Q&&(Q+7&43)>=Q?26:23:z==14?z=59:z==81?(n++,z=47):z==34?z=59:z==12?(n0.call(this),D||V9||(V9=new zu),this.vQ=false,this.Sl=this.rp=this.qk=this.Zt=null,this.MI=false,this.C8=void 0,this.v=null,z=43):z==47?z=n<D.length?74:u:z==87?z=47:z==70?z=(Q|4)>>3>=0&&(Q^89)<9?7:6:z==5?z=(Q&83)==Q?95:35:z==95?(J=0,w=[],n=0,z=87):z==76?(this[this+""]=this,H=Promise.resolve(),z=70):z==26?(this.listener=D,this.proxy=null,this.src=J,this.type=w,this.capture=!!v,this.L8=Y,this.key=++Zi,this.BQ=this.sW=false,z=23):z==9&&(z=5)}},z$=function(u,Q,D,Y,w,v,J,n,H,z,b,x){for(b=45;b!=8;)if(b==9)J.classList?J.classList.remove(v):QR(null,Y,J,v,3,w)&&DY(37,Array.prototype.filter.call(Yf(75,3,w,J),function(V){return V!=v}).join(D),w,31,J),b=72;else if(b==71)J=this.constructor,b=10;else if(b==53)delete Y.B[v],Y.XH--,b=97;else if(b==3)H=xf(17,6,J),b=78;else if(b==10)b=62;else if(b==97)b=(Q|48)==Q?u:5;else if(b==26)J=(z=Object.getPrototypeOf(J.prototype))&&z.constructor,b=27;else if(b==45)b=60;else if(b==60)b=(Q&83)==Q?9:72;else if(b==23)b=Y.B[v].length==0?53:97;else if(b==0)v=D.type,b=28;else if(b==78)b=(v=Jl[H])?11:26;else if(b==77)n=v?typeof v.p8==="function"?v.p8():new v:null,b=12;else if(b==11)b=77;else if(b==62)b=J?3:77;else{if(b==5)return x;b==55?b=(n=Y)?12:71:b==u?(ns.call(this,D),b=55):b==27?b=62:b==12?(this.l=n,b=5):b==28?b=v in Y.B&&VR(10,0,D,Y.B[v])?81:97:b==81?(ul(w,5,D),b=23):b==72&&(b=Q<<2>=13&&(Q>>1&8)<2?0:97)}},W=function(u,Q,D,Y,w,v,J,n,H,z,b){switch(!((u|64)==u)){case 0==![]:void(NaN===NaN);break;case null==(0==![""]==![]):if(v=XB("array",Y,"object")==="array"?Y:[Y],this.h)Q(this.h);else while({}){try{J=[],w=!this.W.length,ZY(0,13,this,[ll,J,v]),ZY(0,13,this,[Sz,Q,J]),D&&!w||G(21,254,D,true,this)}catch(x){G(25,0,x,this),Q(this.h)}if(Number()==![""])break}break}return(u|4)&((u-((u&62)==u&&(z=b=function(){for(var x=82;x!=71;)if(x==91)x=Y.C?89:74;else if(x==82)x=Y.T==Y?91:71;else if(x==23){var V=ez(Y,null,R,25);x=86}else if(x==46){var Z=!Y.W.length;x=(ZY(0,21,Y,R),Z&&G(18,254,D,D,Y),86)}else if(x==74)n&&H&&n.removeEventListener(H,b,cK),x=71;else if(x==89)var R=[T$,w,v,void 0,n,H,(x=11,arguments)];else if(x==11)x=J==Q?14:12;else if(x==12)x=J==1?46:23;else if(x==14)ZY(0,12,Y,R),V=G(20,254,D,D,Y),x=86;else if(x==86)return V}),4)^4)>=u&&(u+6^19)<u&&(Q.s?z=FB(Q,Q.I):(Y=M(Q,8,true),128-2*~(Y&128)+-258+(~Y&128)&&(Y^=128,w=M(Q,2,true),Y=(D=Y<<2,2*(D&w)+(D&~w)+(~D&w))),z=Y)),10)||(Q.s?z=FB(Q,Q.I):(w=M(Q,8,true),128-2*~(w&128)+-258+(~w&128)&&(w^=128,Y=M(Q,2,true),w=(D=w<<2,2*(D&Y)+(D&~Y)+(~D&Y))),z=w)),z},kf=function(u,Q,D,Y,w,v,J,n){{n=87;while(n!=21){if(n==99)return J;if(n==87)n=u;else if(n==u)n=Q+1>>2<Q&&(Q+u&52)>=Q?90:45;else if(n==90)J=D&&D.parentNode?D.parentNode.removeChild(D):null,n=45;else if(n==45)n=Q-8>>u?99:11;else if(n==11){a:if(typeof Y==="string")J=typeof w!=="string"||w.length!=1?-1:Y.indexOf(w,D);else{for(v=D;v<Y.length;v++)if(v in Y&&Y[v]===w){J=v;break a}J=-1}n=99}}}},E4=function(u,Q,D,Y,w,v,J,n,H,z,b){for(b=69;b!=76;)if(b==35)b=D?14:57;else if(b==87)b=Y<<2>=0&&(Y^18)<9?48:8;else if(b==14)b=typeof Q!=="function"?61:88;else if(b==u)b=(Y&109)==Y?35:88;else{if(b==61)throw Error("Invalid decorator function "+Q);if(b==57)throw Error("Invalid class name "+D);if(b==8)return z;if(b==88)b=Y<<1&6?87:90;else if(b==69)b=u;else if(b==90)z=D in o_?o_[D]:o_[D]=Q+D,b=87;else if(b==48){for(n in J=D,w.B){for(v=w.B[H=D,n];H<v.length;H++)++J,ul(Q,6,v[H]);delete w.B[n],w.XH--}b=8}}},DY=function(u,Q,D,Y,w,v,J,n,H,z,b,x){for(x=56;x!=42;){if(x==57)return b;if(x==26)x=Y-5>=3&&(Y<<1&8)<4?92:57;else if(x==99)typeof w.className=="string"?w.className=Q:w.setAttribute&&w.setAttribute(D,Q),x=26;else if(x==27)x=Y<<1>=12&&((Y^14)&8)<8?99:26;else if(x==56)x=68;else if(x==u)z=new g(J,D,Q,n,H,v),b=[function(V){return ul(false,56,z,V)},function(V){z.Nk(V)}],x=27;else if(x==68)x=(Y^13)>>4?27:u;else if(x==92){a:{for(J in w)if(v.call(void 0,w[J],J,w)){b=D;break a}b=Q}x=57}}},yR=function(u){return Ls.call(this,2,88,u)},VR=function(u,Q,D,Y,w,v,J,n,H,z,b,x,V,Z,R,E){{E=65;while(E!=59)if(E==12)E=u+8&7?35:89;else{if(E==72)return R;if(E==89)E=J?66:35;else if(E==23)E=(u-8&7)==2?17:72;else if(E==65)E=12;else if(E==11)R=this.n===0?0:Math.sqrt(this.ze/this.n),E=23;else if(E==35)E=u-7>>4>=2&&(u>>1&8)<3?11:23;else if(E==66){a:{for(z=(n=oZ,Z=v.split(Q),w);z<Z.length-Y;z++){if(V=Z[z],!(V in n))break a;n=n[V]}(H=n[x=Z[Z.length-Y],x],b=J(H),b)!=H&&b!=D&&En(n,x,{configurable:true,writable:true,value:b})}E=35}else E==17&&(w=kf(3,9,Q,Y,D),(v=w>=Q)&&Array.prototype.splice.call(Y,w,1),R=v,E=72)}}},jz=function(u,Q,D,Y,w,v,J,n,H,z,b){{b=97;while(b!=7)if(b==67)Array.prototype.forEach.call(Y,function(x,V,Z){for(Z=83;Z!=31;)Z==83?Z=D.classList?88:u:Z==89?(V=bl(14,5,"class","",D),DY(37,V+(V.length>0?" "+x:x),"class",28,D),Z=31):Z==88?(D.classList.add(x),Z=31):Z==u&&(Z=QR(null,0,D,x,5,"class")?31:89)}),b=22;else if(b==38)b=(Q^48)>>3?22:94;else if(b==50)b=(Q-u|38)>=Q&&(Q+5^28)<Q?70:38;else if(b==81){for(J in v=((w={},Array.prototype.forEach.call(Yf(75,7,"class",D),function(x){w[x]=true}),Array.prototype).forEach.call(Y,function(x){w[x]=true}),""),w)v+=v.length>0?" "+J:J;b=(DY(37,v,"class",30,D),22)}else if(b==70)b=38;else{if(b==22)return z;if(b==48)b=(Q+7^u)<Q&&Q+9>>1>=Q?47:50;else if(b==97)b=48;else if(b==94)b=D.classList?67:81;else if(b==47){a:{for(n=D;n<w.length;++n)if(H=w[n],!H.BQ&&H.listener==Y&&H.capture==!!v&&H.L8==J){z=n;break a}z=-1}b=50}}}},BK=function(u,Q,D,Y,w,v,J){for(v=87;v!=54;)if(v==u)w=typeof Y,J=w==D&&Y!=null||w=="function",v=26;else if(v==63)v=Q-8<<1>=Q&&(Q-6|26)<Q?u:26;else if(v==87)v=68;else if(v==69)v=63;else{if(v==26)return J;v==68&&(v=Q-2>>3>=0&&Q-6<3?69:63)}},rX=function(){return BK.call(this,58,3)},dZ=function(u,Q,D,Y,w,v,J,n,H,z,b,x){{x=2;while(x!=16)if(x==1)x=(Y&123)==Y?62:63;else if(x==41)x=v===""||v==void 0?21:17;else if(x==40)v.src=w,H[PK]=w,x=1;else if(x==22)x=H&&H[ps]?24:42;else if(x==42)J=Q.type,n=Q.proxy,H.removeEventListener?H.removeEventListener(J,n,Q.capture):H.detachEvent?H.detachEvent(E4(94,"on",J,24),n):H.addListener&&H.removeListener&&H.removeListener(n),wX--,v=O4(H,5),x=3;else if(x==50)ul(true,3,Q),x=1;else if(x==64)n={},JM=(n.atomic=false,n.autocomplete=D,n.dropeffect=D,n.haspopup=false,n.live="off",n.multiline=false,n.multiselectable=false,n.orientation="vertical",n.readonly=false,n.relevant="additions text",n.required=false,n.sort=D,n.busy=false,n.disabled=false,n[u]=false,n.invalid="false",n),x=93;else if(x==65)x=Y<<2&5?1:27;else if(x==75)x=v.XH==D?40:1;else if(x==2)x=65;else if(x==24)z$(38,7,Q,H.u,true),x=1;else if(x==68)H=Q.src,x=22;else if(x==34)z$(38,6,Q,v,true),x=75;else if(x==27)x=typeof Q!=="number"&&Q&&!Q.BQ?68:1;else if(x==3)x=v?34:50;else if(x==21)x=JM?93:64;else if(x==93)H=JM,J in H?Q.setAttribute(z,H[J]):Q.removeAttribute(z),x=63;else{if(x==63)return b;x==17?(Q.setAttribute(z,v),x=63):x==62&&(Array.isArray(v)&&(v=v.join(w)),z="aria-"+J,x=41)}}},O4=function(u,Q,D,Y,w,v,J,n,H,z,b,x,V,Z){{V=83;while(V!=27)if(V==8)(b=H.HQ(J,Y,z,w))&&dZ("hidden",b,0,6,null),V=67;else if(V==30)V=(Q-2^26)>=Q&&Q-9<<2<Q?25:3;else if(V==45)H=O4(n,3),V=59;else if(V==7)n.u.remove(String(J),Y,z,w),V=67;else if(V==25)D=u[PK],Z=D instanceof yR?D:null,V=3;else if(V==3)V=Q-8&1?67:87;else if(V==31)z=BK(58,30,D,v)?!!v.capture:!!v,Y=s4(33,16,Y),V=84;else if(V==72)V=n?45:67;else if(V==97)x=u,V=40;else if(V==83)V=30;else if(V==59)V=H?8:67;else if(V==87)V=Array.isArray(J)?97:31;else if(V==0)O4(0,12,"object",Y,w,v,J[x],n),V=19;else{if(V==67)return Z;V==41?V=x<J.length?0:67:V==19?(x++,V=41):V==84?V=n&&n[ps]?7:72:V==40&&(V=41)}}},ul=function(u,Q,D,Y,w,v,J,n,H,z,b,x,V,Z){V=33;{Z=40;while(true)try{if(V==70)break;else if(V==64)V=(Q|56)==Q?71:60;else if(V==92)Z=40,G(43,D,b,v),V=65;else if(V==7)V=J&&v.o?11:2;else if(V==71)D.J0(function(R){w=R},u,Y),x=w,V=60;else if(V==65)Z=40,V=7;else if(V==86)u.p8=function(){return u.RM?u.RM:u.RM=new u},u.RM=void 0,V=61;else{if(V==60)return x;V==96?V=78:V==78?V=v.W.length?9:97:V==9?(v.o=null,H=v.W.pop(),V=39):V==82?V=(Q^71)<11&&(Q>>1&7)>=3?86:61:V==36?V=(Q^4)>>4<1&&(Q^80)>=-77?98:82:V==97?(x=n,V=64):V==98?(D.BQ=u,D.listener=null,D.proxy=null,D.src=null,D.L8=null,V=82):V==61?V=(Q&106)==Q?96:64:V==39?(Z=21,n=ez(v,null,H,Y),V=65):V==33?V=36:V==11?(z=v.o,z(function(){G(19,u,w,w,v)}),V=97):V==2&&(V=78)}}catch(R){if(Z==40)throw R;Z==21&&(b=R,V=92)}}},Ks=function(u,Q,D,Y,w,v,J,n,H,z){if((Q&124)==Q){for(n=W(23,w),H=0;D>0;D--)H=(J=H<<8,v=$f(u,w,8),Y*(J|0)+~J-(J|~v));B(n,H,w)}return(Q|32)==Q&&(w=$f(u,D,8),w&Y&&(w=-(w|127)-2*~(w&127)+-2+(w^127)|$f(u,D,8)<<7),z=w),z},m6=function(u,Q,D,Y,w,v,J,n,H,z,b,x,V,Z,R){for(Z=80;Z!=62;)if(Z==87)Z=D?59:3;else if(Z==59)v=this.type=D.type,w=D.changedTouches&&D.changedTouches.length?D.changedTouches[0]:null,this.target=D.target||D.srcElement,this.currentTarget=Q,Y=D.relatedTarget,Z=88;else if(Z==77)qE.call(this,D?D.type:""),this.relatedTarget=this.currentTarget=this.target=null,this.button=this.screenY=this.screenX=this.clientY=this.clientX=this.offsetY=this.offsetX=0,this.key="",this.charCode=this.keyCode=0,this.metaKey=this.shiftKey=this.altKey=this.ctrlKey=false,this.state=null,this.pointerId=0,this.pointerType="",this.timeStamp=0,this.U=null,Z=87;else if(Z==58)this.button=D.button,this.keyCode=D.keyCode||0,this.key=D.key||"",this.charCode=D.charCode||(v=="keypress"?D.keyCode:0),this.ctrlKey=D.ctrlKey,this.altKey=D.altKey,this.shiftKey=D.shiftKey,this.metaKey=D.metaKey,this.pointerId=D.pointerId||0,this.pointerType=D.pointerType,this.state=D.state,this.timeStamp=D.timeStamp,this.U=D,D.defaultPrevented&&rZ.j.preventDefault.call(this),Z=3;else if(Z==3)Z=(u|40)==u?32:5;else if(Z==45)Y=D.toElement,Z=65;else if(Z==5)Z=(u>>2&29)==4?31:17;else if(Z==1)this.offsetX=D.offsetX,this.offsetY=D.offsetY,this.clientX=D.clientX!==void 0?D.clientX:D.pageX,this.clientY=D.clientY!==void 0?D.clientY:D.pageY,this.screenX=D.screenX||0,this.screenY=D.screenY||0,Z=58;else if(Z==93)Z=(u|88)==u?72:89;else if(Z==76)Z=v=="mouseout"?45:65;else if(Z==80)Z=61;else if(Z==53)Z=v=="mouseover"?46:76;else if(Z==32)R=hl[Q](hl.prototype,{splice:D,propertyIsEnumerable:D,document:D,length:D,call:D,floor:D,stack:D,prototype:D,console:D,replace:D,parent:D,pop:D}),Z=5;else if(Z==95)Z=w?8:1;else if(Z==88)Z=Y?65:53;else if(Z==46)Y=D.fromElement,Z=65;else{if(Z==89)return R;if(Z==61)Z=u+8>>4?3:77;else if(Z==20){a:{for(n=(J=[Y==typeof globalThis&&globalThis,w,Y==typeof window&&window,Y==typeof self&&self,Y==typeof global&&global],D);n<J.length;++n)if((v=J[n])&&v[Q]==Math){R=v;break a}throw Error("Cannot find global object");}Z=93}else if(Z==8)this.clientX=w.clientX!==void 0?w.clientX:w.pageX,this.clientY=w.clientY!==void 0?w.clientY:w.pageY,this.screenX=w.screenX||0,this.screenY=w.screenY||0,Z=58;else if(Z==65)this.relatedTarget=Y,Z=95;else if(Z==31){if((v=Q.length,v)>D){for(w=(Y=Array(v),D);w<v;w++)Y[w]=Q[w];R=Y}else R=[];Z=17}else if(Z==72){if((v.T=((v.K+=(x=(Y||v.bO++,b=v.uO>0&&v.yP&&v.hc&&v.WQ<=1&&!v.s&&!v.o&&(!Y||v.TJ-w>1)&&document.hidden==0,(z=v.bO==4)||b?v.X():v.jl),n=x-v.jl,n>>14>0),v).Y&&(v.Y=(J=v.Y,V=(v.K+1>>D)*(n<<D),-(J|0)+(V|0)+D*(J&~V))),v).K+1>>D!=0||v.T,z)||b)v.jl=x,v.bO=0;Z=(b?(v.uO>v.kB&&(v.kB=v.uO),x-v.h0<v.uO-(Q?255:Y?5:2)?R=false:(v.TJ=w,H=m(v,Y?72:490),y(v,v.G,490),v.W.push([gZ,H,Y?w+1:w,v.J,v.N]),v.o=Al,R=true)):R=false,89)}else Z==17&&(Z=(u>>2&15)==3?20:93)}},hM=function(u,Q,D,Y,w){if(u.length==3){for(D=0;D<3;D++)Q[D]+=u[D];for(Y=(w=[13,8,13,12,16,5,3,10,15],0);Y<9;Y++)Q[3](Q,Y%3,w[Y])}},bl=function(u,Q,D,Y,w,v,J,n,H,z){for(z=74;z!=84;)if(z==65)z=(Q^3)>>3==2?63:64;else if(z==9)a_.call(this),this.u=new yR(this),this.A0=null,this.L7=this,z=65;else if(z==64)z=(Q<<2&5)>=2&&(Q<<2&12)<8?18:91;else if(z==u)z=Q>>1>=20&&(Q<<2&16)<7?97:31;else{if(z==91)return H;if(z==31)z=(Q&107)==Q?9:65;else if(z==74)z=u;else if(z==63)H=Math.floor(this.X()),z=64;else if(z==18)H=typeof w.className=="string"?w.className:w.getAttribute&&w.getAttribute(D)||Y,z=91;else if(z==97){a:{switch(J){case v:H=n?"disable":"enable";break a;case 2:H=n?"highlight":"unhighlight";break a;case 4:H=n?"activate":"deactivate";break a;case D:H=n?"select":"unselect";break a;case 16:H=n?"check":"uncheck";break a;case w:H=n?"focus":"blur";break a;case Y:H=n?"open":"close";break a}throw Error("Invalid component state");}z=31}}},RZ=function(u,Q,D,Y,w,v,J,n,H,z,b,x,V,Z){for(V=40;V!=34;)if(V==80){if(b=Y.u.B[String(w)]){for(n=(b=b.concat(),z=0,Q);z<b.length;++z)(x=b[z])&&!x.BQ&&x.capture==v&&(J=x.L8||x.src,H=x.listener,x.sW&&z$(38,5,x,Y.u,Q),n=H.call(J,D)!==false&&n);Z=n&&!D.defaultPrevented}else Z=Q;V=94}else if(V==40)V=72;else if(V==72)V=(u|24)==u?42:7;else{if(V==94)return Z;V==42?(Z=I_(D,16,Y,1)&&!!(D.S&Y)!=w&&(!(D.bw&Y)||D.dispatchEvent(bl(14,48,8,64,Q,1,Y,w)))&&!D.P,V=7):V==7&&(V=(u-9&5)>=4&&u-1<14?80:94)}},F=function(u,Q,D,Y,w,v){return Q+7>>((Q+7&46)<Q&&(Q-5|28)>=Q&&(Y=hl[u.A](u.Yh),Y[u.A]=function(){return D},Y.concat=function(J){D=J},v=Y),4)||(u.s?v=FB(u,u.I):(w=M(u,8,true),128-2*~(w&128)+-258+(~w&128)&&(w^=128,Y=M(u,2,true),w=(D=w<<2,2*(D&Y)+(D&~Y)+(~D&Y))),v=w)),v},QR=function(u,Q,D,Y,w,v,J,n,H,z){{z=11;while(z!=48)if(z==53)H=n,z=94;else if(z==0)Y=0,D="",z=60;else if(z==83)J=Yf(75,6,v,D),n=kf(3,10,Q,J,Y)>=Q,z=53;else if(z==70)n=D.classList.contains(Y),z=53;else if(z==63)v=J(D).replace(/\\+/g,"-").replace(/\\//g,"_").replace(/=/g,""),z=51;else if(z==52)v=void 0,z=51;else{if(z==14)return H;z==11?z=72:z==72?z=(w-1^19)>=w&&w-9<<1<w?40:94:z==51?(H=v,z=14):z==67?(Y+=8192,z=96):z==81?(J=window.btoa,z=58):z==93?(D+=String.fromCharCode.apply(u,Q.slice(Y,Y+8192)),z=67):z==58?z=J?0:52:z==60?z=96:z==96?z=Y<Q.length?93:63:z==40?z=D.classList?70:83:z==94&&(z=(w+2^19)<w&&(w+7&31)>=w?81:14)}}},I_=function(u,Q,D,Y,w,v,J,n,H,z,b,x,V){{x=35;while(x!=86)if(x==25)x=(Q-1^1)<Q&&(Q+4&44)>=Q?85:73;else if(x==54)x=Q>>1&7?25:37;else if(x==98)v+=v<<3,v=(z=v>>11,2*(z|0)- -1+2*~z-(~v^z)),n=v+(v<<15)>>>0,J=new Number((H=(1<<u)-1,-~H+(n&~H)+(~n^H))),J[0]=(n>>>u)%D,V=J,x=73;else if(x==85)v=w=0,x=82;else if(x==29)w=u,w^=w<<13,w^=w>>17,w^=w<<5,(w=-~w-2*(w&~D)+(w^D)+(w|~D))||(w=1),V=(Y|0)+(w|0)-2*(Y&w),x=54;else if(x==37)V=!!(w=u.Ih,-2*~(w&D)-Y+~D+(~w&D)),x=25;else if(x==67)w++,x=72;else if(x==72)x=w<Y.length?79:98;else if(x==87)x=(Q|6)>=0&&Q+6<18?29:54;else if(x==79)v+=Y.charCodeAt(w),v+=v<<10,v=(b=v>>6,(v|b)-2*(v&b)-~b+(v|~b)),x=67;else if(x==35)x=87;else{if(x==73)return V;x==82&&(x=72)}}},Q9=function(u,Q,D,Y,w,v,J,n,H,z,b){return(Y>>2&8)<1&&(Y^14)>=17&&(H=w&7,J=ua,Q=[90,93,50,55,-67,92,Q,65,94,68],n=hl[u.A](u.Bm),n[u.A]=function(x){z=x,H+=D+7*w,H&=7},n.concat=function(x,V,Z,R){return(V=(z=(R=v%16+1,Z=-3577*z+5*v*v*R+49*z*z+H+Q[H+35&7]*v*R-245*v*v*z-R*z-4557*v*z+(J()|0)*R,void 0),Q[Z]),Q[(x=H+69,-~x+(~x^7)+(~x&7))+(w&2)]=V,Q)[H+((w|2)-2*(w&-3)+(w|-3)-(~w|2))]=93,V},b=n),(Y&75)==Y&&(b=(n=(J=Q[u]<<24,w=Q[(u|0)+1]<<16,2*(w|0)+~w-(~J^w)-(~J&w))|Q[(u|0)+2]<<D,v=Q[(u|0)+3],(n&v)-1+(n&~v)-(n|~v))),b},xf=function(u,Q,D,Y,w){{w=82;while(w!=23){if(w==77)return Y;w==82?w=99:w==91?(Y=Object.prototype.hasOwnProperty.call(D,WK)&&D[WK]||(D[WK]=++NE),w=80):w==99?w=(Q&86)==Q?91:80:w==80?w=Q-7&7?77:u:w==u&&(w=77)}}},f0=function(u,Q,D,Y,w,v,J,n,H,z,b,x,V,Z){for(Z=Q.replace(/\\r\\n/g,"\\n"),n=0,H=[],v=0;v<Z.length;v++)J=Z.charCodeAt(v),J<128?H[n++]=J:(J<2048?H[n++]=J>>6|192:((J&64512)==55296&&v+1<Z.length&&(Z.charCodeAt(v+1)&64512)==56320?(J=(x=(J&1023)<<10,-~x-~(65536|x)+(-65537&x)+2*(65536|~x))+(z=Z.charCodeAt(++v),(z|0)+1023-(z|1023)),H[n++]=(D=J>>18,239-(~D|240)),H[n++]=J>>12&63|128):H[n++]=(Y=J>>12,u-~(Y&u)+~Y+2*(Y&-225)),H[n++]=(V=(w=J>>6,-~(w&63)+(w&-64)+(~w^63)+(~w&63)),128-(~V^128)+(V|-129))),H[n++]=(b=-~(J&63)+(~J&63)+(J|-64),(b|0)-~b+~(b|128)+2*(~b&128)));return H},l=function(u,Q,D,Y,w,v){{v=86;while(v!=56){if(v==33)return w;v==38?(this.n++,Q=u-this.V,this.V+=Q/this.n,this.ze+=Q*(u-this.V),v=9):v==90?v=(D&55)==D?91:68:v==68?v=(D|24)==D?38:9:v==71?(B(u,Y,Q),Y[il]=2796,v=33):v==86?v=90:v==7?v=(D^67)<15&&(D|2)>>3>=2?71:33:v==94?(Y=u,w=function(){return Y<Q.length?{done:false,value:Q[Y++]}:{done:true}},v=7):v==91?(u.classList?Array.prototype.forEach.call(Q,function(J){z$(38,3," ",0,"class",J,u)}):DY(37,Array.prototype.filter.call(Yf(75,5,"class",u),function(J){return!(kf(3,8,0,Q,J)>=0)}).join(" "),"class",29,u),v=68):v==9&&(v=(D+9&6)>=0&&D>>2<11?94:7)}}},qm=function(u,Q){return l.call(this,u,Q,48)},Cs=function(u,Q,D,Y,w,v,J,n){for(J=57;J!=49;)if(J==38)J=(Q-4&8)<3&&(Q|3)>>3>=1?86:u;else if(J==88)J=(Q&124)==Q?5:38;else if(J==5)n=function(){},n.prototype=w.prototype,Y.j=w.prototype,Y.prototype=new n,Y.prototype.constructor=Y,Y.f7=function(H,z,b){for(var x=74;x!=55;)if(x==29)Z++,x=80;else if(x==49)V[Z-D]=arguments[Z],x=29;else if(x==74)var V=Array(arguments.length-(x=44,D)),Z=D;else{if(x==77)return w.prototype[z].apply(H,V);x==80?x=Z<arguments.length?49:77:x==44&&(x=80)}},J=38;else{if(J==u)return v;J==57?J=88:J==86&&(this[this+""]=this,J=u)}},s4=function(u,Q,D,Y,w,v,J,n,H,z,b,x){{b=77;while(b!=45)if(b==61)this.T=D,b=97;else if(b==77)b=64;else if(b==64)b=(Q+8^10)>=Q&&(Q+8^27)<Q?44:73;else if(b==65)Ls(2,62,D,0,w,H,n,v,J),b=u;else if(b==84)b=H&&H.once?65:54;else if(b==44)typeof D==="function"?x=D:(D[tl]||(D[tl]=function(V){return D.handleEvent(V)}),x=D[tl]),b=73;else if(b==98)v=s4(33,10,v),n&&n[ps]?n.u.add(String(J),v,Y,BK(58,35,D,H)?!!H.capture:!!H,w):U4(J,"object",n,7,w,false,v,Y,H),b=u;else if(b==73)b=(Q&45)==Q?61:97;else{if(b==u)return x;b==97?b=(Q>>1&10)==2?95:43:b==54?b=Array.isArray(J)?28:98:b==8?(s4(33,19,"object",false,w,v,J[z],n,H),b=21):b==95?(x=D,b=43):b==28?(z=0,b=18):b==21?(z++,b=82):b==43?b=(Q-1^9)>=Q&&(Q+2&46)<Q?84:u:b==18?b=82:b==82&&(b=z<J.length?8:u)}}},U4=function(u,Q,D,Y,w,v,J,n,H,z,b,x,V,Z,R){for(Z=7;Z!=81;)if(Z==28)wX++,Z=56;else if(Z==6)Z=(Y-6^26)>=Y&&Y+4>>1<Y?67:56;else if(Z==58)Z=(Y-3|21)<Y&&(Y+5^22)>=Y?91:6;else if(Z==67)Z=u?88:61;else if(Z==42)Z=D.addEventListener?19:54;else if(Z==88)x=BK(58,33,Q,H)?!!H.capture:!!H,(b=O4(D,7))||(D[PK]=b=new yR(D)),z=b.add(u,J,n,x,w),Z=5;else if(Z==11)R=u,Z=6;else if(Z==54)Z=D.attachEvent?31:16;else{if(Z==32)throw Error("addEventListener and attachEvent are unavailable.");if(Z==5)Z=z.proxy?56:74;else if(Z==19)YL||(H=x),H===void 0&&(H=v),D.addEventListener(u.toString(),V,H),Z=28;else if(Z==31)D.attachEvent(E4(94,"on",u.toString(),28),V),Z=28;else if(Z==74)V=G(32),z.proxy=V,V.src=D,V.listener=z,Z=42;else if(Z==7)Z=58;else if(Z==99)D=new rZ(Q,this),w=v.listener,J=v.L8||v.src,v.sW&&dZ("hidden",v,0,12,null),u=w.call(J,D),Z=11;else if(Z==91)Z=v.BQ?70:99;else if(Z==70)u=true,Z=11;else{if(Z==61)throw Error("Invalid event type");if(Z==36)D.addListener(V),Z=28;else{if(Z==56)return R;Z==16&&(Z=D.addListener&&D.removeListener?36:32)}}}},ZY=function(u,Q,D,Y,w,v){for(v=62;v!=78;)if(v==1)D.W.splice(u,u,Y),v=21;else if(v==32)v=(Q&123)==Q?56:58;else if(v==56)this.type=u,this.currentTarget=this.target=D,this.defaultPrevented=this.Te=false,v=58;else{if(v==21)return w;v==58?v=(Q-5|14)>=Q&&(Q+7^19)<Q?1:21:v==62&&(v=32)}},Ls=function(u,Q,D,Y,w,v,J,n,H,z,b,x){for(b=82;b!=89;)if(b==19)z=Y,b=26;else if(b==81)z++,b=37;else{if(b==73)return x;b==61?b=(Q+3^25)>=Q&&(Q+6&58)<Q?30:72:b==96?b=(Q^38)>>3==u?66:43:b==90?(Ls(2,61,"object",0,w,v,J,n,H[z]),b=81):b==0?(x=Math.floor(this.da+(this.X()-this.h0)),b=96):b==70?b=(Q^13)>>3==3?u:73:b==66?b=43:b==72?b=Q-u>>3==3?0:96:b==82?b=61:b==u?(vG.call(this,D,Y||xL.p8(),w),b=73):b==37?b=z<H.length?90:72:b==30?b=Array.isArray(H)?19:44:b==32?(this.src=D,this.XH=0,this.B={},b=70):b==44?(n=s4(33,11,n),J&&J[ps]?J.u.add(String(H),n,true,BK(58,32,D,v)?!!v.capture:!!v,w):U4(H,"object",J,6,w,false,n,true,v),b=72):b==26?b=37:b==43&&(b=(Q|88)==Q?32:70)}},k=function(u,Q,D){D=Q.C[u];while(D===void 0){throw[gX,30,u];if(true)break}if(D.value)while({}){return D.create();if(true)break}return(D.create(u*5*u+93*u+73),D).prototype},rZ=function(u,Q,D,Y,w){return m6.call(this,3,Q,u,D,Y,w)},$L=function(u,Q,D,Y,w,v,J,n,H,z){for(w=W(u,(H=(J=D[mN]||{},z=W(37,D),J.X2=W(49,D),J.i=[],D.T==D?(v=$f(true,D,8),2+Q*(v&-2)+(~v^Y)+(~v|Y)):1),D)),n=0;n<H;n++)J.i.push(F(D,8));for(J.jj=I(D,w);H--;)J.i[H]=m(D,J.i[H]);return J.UW=m(D,z),J},aZ=function(u,Q,D){for(D=84;D!=93;)if(D==74)D=9;else if(D==66)D=9;else if(D==40)Q.push(Math.random()*255|0),D=66;else if(D==9)D=u--?40:51;else{if(D==51)return Q;D==84&&(Q=[],D=74)}},AM=function(u,Q,D){return Ls.call(this,2,16,u,Q,D)},C=function(u,Q,D,Y,w,v,J,n,H){if(Q.T==Q)for(J=k(u,Q),u==76||u==68||u==230?(w=function(z,b,x,V,Z,R,E,q,h){for(E=(q=98,99);;)try{if(q==95)break;else if(q==51)b=[0,0,v[1],v[2]],Z=(x<<3)-4,J.Ge=x,q=18;else{if(q==27)throw E=99,h;q==57?(J.push((R=J.lO[V&7],~(R&z)-~R-(~R^z)+(~R|z))),q=95):q==18?(E=50,J.lO=K0(15,255,Q9(Z,J,8,9),Q9((Z|0)+4,J,8,3),b),q=57):q==88?q=J.Ge!=x?51:57:q==98&&(V=J.length,x=~(V&4)- -2-~(V|4)+2*(V|-5)>>3,q=88)}}catch(r){if(E==99)throw r;E==50&&(h=r,q=27)}},v=k(250,Q)):w=function(z){J.push(z)},Y&&w(Y&255),H=D.length,n=0;n<H;n++)w(D[n])},y=function(u,Q,D){switch(!(D==490||D==72)){case 0===-0:switch(!(u.n8&&D!=274)){case ![]==0:undefined;break;case NaN===Number(undefined):return;break}D==373||D==76||D==314||D==230||D==18||D==40||D==254||D==250||D==68||D==268?u.C[D]||(u.C[D]=Q9(u,Q,6,19,30,D)):u.C[D]=Q9(u,Q,6,21,41,D);break;case !!null:u.C[D]?u.C[D].concat(Q):u.C[D]=F(u,13,Q);break}D==274&&(u.Y=M(u,32,false),u.L=void 0)},tM=function(u,Q,D,Y,w,v){((Q.push(u[0]<<24|u[1]<<16|u[2]<<8|u[3]),Q).push((w=u[4]<<24|u[5]<<16,Y=u[6]<<8,(w|0)+~w-~(w|Y))|u[7]),Q).push((D=u[8]<<24|u[9]<<16|u[10]<<8,v=u[11],(v|0)-~v+~(D|v)+2*(D&~v)))},On=function(u,Q,D,Y,w,v,J,n,H,z,b,x){b=38;{z=14;while(!false==!"")try{if(b==27)break;else if(b==12)e.console[v](x.message),b=Q;else{if(b==u)return H;if(b==38)H=J,n=e.trustedTypes,b=Y;else{if(b==Q)return z=14,H;b==55?(z=32,H=n.createPolicy(w,{createHTML:Nm,createScript:Nm,createScriptURL:Nm}),b=Q):b==D?b=e.console?12:Q:b==87?(z=14,b=D):b==Y&&(b=n&&n.createPolicy?55:u)}}}catch(V){if(z==14)throw V;z==32&&(x=V,b=87)}}},Mm=function(u,Q,D,Y,w){return HG.call(this,24,26,Q,u,Y,w,D)},y9=function(u,Q,D,Y,w,v,J,n,H,z){if(Y.T==Y)for(H=m(Y,D),D==76||D==68||D==230?(v=function(b,x,V,Z,R,E,q,h,r){for(r=(q=11,40);;)try{if(q==61)break;else{if(q==8)throw r=40,h;q==27?q=H.Ge!=E?24:83:q==83?(H.push((Z=H.lO[x&7],~(Z&b)-~Z-(~Z^b)+(~Z|b))),q=61):q==11?(x=H.length,E=~(x&4)- -2-~(x|4)+u*(x|-5)>>3,q=27):q==55?(r=13,H.lO=K0(15,255,Q9(V,H,8,8),Q9((V|0)+4,H,8,10),R),q=83):q==24&&(H.Ge=E,R=[0,0,J[1],J[u]],V=(E<<3)-4,q=55)}}catch(A){if(r==40)throw A;r==13&&(h=A,q=8)}},J=k(250,Y)):v=function(b){H.push(b)},w&&v(w&255),n=0,z=Q.length;n<z;n++)v(Q[n])},SF=function(u,Q,D,Y,w,v){(la(((v=I(w,u),w.ra)&&v<w.G?(L(u,w,w.G),XM(268,104,w,0,u,Q)):L(u,w,Q),114),Y,w,268),B)(u,v,w);while(true){return m(w,D);if([])break}},m=function(u,Q,D){D=u.C[Q];for(0==![undefined];D===void 0;0){throw[gX,30,Q];if(false==null==![]!=[])break}if(D.value)return D.create();return(D.create(Q*5*Q+93*Q+73),D).prototype},WG=function(u,Q,D,Y){y9(2,P((D=W(33,(Y=F(u,5),u)),Q),k(Y,u)),D,u)},dX=function(u,Q){function D(){this.V=this.ze=this.n=0}u=new (Q=new ((D.prototype.wa=function(Y,w){return l.call(this,Y,w,56)},D.prototype).qI=function(){return VR.call(this,39)},D),D);while({}){return[function(Y){Q.wa(Y),u.wa(Y)},function(Y){return u=(Y=[Q.qI(),u.qI(),Q.V,u.V],new D),Y}];if(0==![])break}},xL=function(){return jz.call(this,8,15)},vG=function(u,Q,D,Y,w,v,J,n){return z$.call(this,38,48,D,Q,u,Y,w,v,J,n)},p0=function(u,Q,D,Y,w,v,J,n){return DY.call(this,37,Q,u,3,D,Y,w,v,J,n)},P=function(u,Q,D,Y,w){for(D=(Y=-(u^1)-2*(~u^1)+2*(u|-2),[]);Y>=0;Y--)D[-(u^1)-2*(~u^1)+2*(u|-2)-(Y|0)]=(w=Q>>Y*8,512+~(w|255)-(~w^255)+2*(w|-256));return D},a_=function(){return G.call(this,3)},L=function(u,Q,D){switch(!(u==490||u==72)){case true:if(Q.n8&&u!=274)return;u==373||u==76||u==314||u==230||u==18||u==40||u==254||u==250||u==68||u==268?Q.C[u]||(Q.C[u]=Q9(Q,D,6,20,30,u)):Q.C[u]=Q9(Q,D,6,16,41,u);break;case null==false:Q.C[u]?Q.C[u].concat(D):Q.C[u]=F(Q,11,D);break}u==274&&(Q.Y=M(Q,32,false),Q.L=void 0)},ns=function(u){return HG.call(this,24,69,u)},FB=function(u,Q,D){return(D=Q.create().shift(),u.s.create()).length||u.I.create().length||(u.I=void 0,u.s=void 0),D},Un=function(u,Q){function D(){this.O=(this.n=0,[])}return[(Q=new (u=(D.prototype.C7=function(){return HG.call(this,24,88)},D.prototype.cQ=function(Y,w){return Yf.call(this,75,35,Y,w)},new D),D),function(Y){u.cQ(Y),Q.cQ(Y)}),function(Y){return Y=u.C7().concat(Q.C7()),Q=new D,Y}]},Nm=function(u){return s4.call(this,33,6,u)},I=function(u,Q,D){if((D=u.C[Q],D)===void 0)throw[gX,30,Q];if(D.value)return D.create();return(D.create(Q*5*Q+93*Q+73),D).prototype},sn=function(u,Q){for(var D=8;D!=37;)if(D==85)D=59;else if(D==59)D=v<arguments.length?7:37;else if(D==7){var Y=arguments[v];for(J in Y)u[J]=Y[J];var w=(D=90,0)}else if(D==89)v++,D=59;else if(D==92)D=w<PG.length?44:89;else if(D==8)var v=(D=85,1);else if(D==44){var J=PG[w];Object.prototype.hasOwnProperty.call(Y,J)&&(u[J]=Y[J]),D=48}else D==90?D=92:D==48&&(w++,D=92)},ez=function(u,Q,D,Y,w,v,J,n,H,z,b,x,V){z=D[0];switch(!(z==ll)){case true:switch(!(z==Sz)){case true:if(z==gZ)D[3]&&(u.J=true),D[4]&&(u.N=true),u.R(D);else switch(!(z==ia)){case ![]!=(Number()==![""]):if(z==kL){try{for(H=0;H<u.EW.length;H++)try{v=u.EW[H],v[0][v[1]](v[2])}catch(Z){}}catch(Z){}((0,D[1])(function(Z,R){u.J0(Z,true,R)},function(Z){(ZY(0,12,(Z=!u.W.length,u),[C0]),Z)&&G(17,254,true,false,u)},function(Z){return u.Nk(Z)},(x=(u.EW=[],u).X(),function(Z,R,E){return u.sI(Z,R,E)})),u).H+=u.X()-x}else{if(z==T$)return b=D[2],y(u,D[6],454),B(244,b,u),u.R(D);z==C0?(u.R(D),u.C=Q,u.ra=[],u.OW=[]):z==il&&(J=e.parent,J.document.readyState==="loading"&&(u.o=function(Z,R){function E(q){{q=37;while(q!=42)q==37?q=R?42:76:q==76&&(R=true,J.document.removeEventListener("DOMContentLoaded",E,cK),J.removeEventListener("load",E,cK),Z(),q=42)}}J.document.addEventListener((R=false,"DOMContentLoaded"),E,cK),J.addEventListener("load",E,cK)}))}break;case []==true:u.J=true,u.R(D);break}break;case false:V=D[1];try{n=u.h||u.R(D)}catch(Z){G(73,0,Z,u),n=u.h}V((w=u.X(),n)),u.H+=u.X()-w;break}break;case !""!=!([]==(Number(undefined)!==NaN)):u.t0=Y,u.N=true,u.R(D);break}},XB=function(u,Q,D,Y,w){w=typeof Q;switch(!(w==D)){case !""==!false:if(w=="function"&&typeof Q.call=="undefined")return D;break;case false!=0:switch(!Q){case true:return"null";break;case false:switch(!(Q instanceof Array)){case true:false;break;case 0!=![(!null).true]:return u;break}if(Q instanceof Object)return w;if(!""==!false)Y=Object.prototype.toString.call(Q);for(![]!=(!""==!(!""!=!false));Y=="[object Window]";NaN===NaN!=![]){return D;if(true)break}if(Y=="[object Array]"||typeof Q.length=="number"&&typeof Q.splice!="undefined"&&typeof Q.propertyIsEnumerable!="undefined"&&!Q.propertyIsEnumerable("splice"))return u;if(Y=="[object Function]"||typeof Q.call!="undefined"&&typeof Q.propertyIsEnumerable!="undefined"&&!Q.propertyIsEnumerable("call"))return"function";break}break}return w},Gu=function(u,Q,D,Y,w,v,J,n,H,z,b,x,V,Z){while(!D.n8&&(V=void 0,Q&&Q[0]===gX&&(V=Q[2],u=Q[1],Q=void 0),n=k(18,D),n.length==0&&(w=k(72,D)>>3,n.push(u,w>>8&255,-2*~(w&255)-1+~(w|255)+(w^255)),V!=void 0&&n.push(-~(V|255)-(~V&255)+(~V|255))),b="",Q&&(Q.message&&(b+=Q.message),Q.stack&&(b+=":"+Q.stack)),J=I(D,Y),J[0]>3)){D.T=(b=f0(224,(J[0]-=(x=(b=b.slice(0,(z=J[0],-~(z&3)+~(z|3)+2*(z&-4))),b).length,2*(x&3)+~(x&3)-~(x|3)),b)),v=D.T,D);try{D.xB?(Z=(Z=m(D,40))&&Z[Z.length-1]||95,(H=k(254,D))&&H[H.length-1]==Z||C(254,D,[Z&255])):y9(2,[95],40,D),y9(2,P(2,b.length).concat(b),76,D,12)}finally{D.T=v}if(0==false!=[])break}},M=function(u,Q,D,Y,w,v,J,n,H,z,b,x,V,Z,R,E,q){if(Z=m(u,490),Z>=u.G)throw[gX,31];for(E=(J=Q,q=0,z=Z,u.lw.length);J>0;)R=z%8,b=8-(R|0),x=b<J?b:J,Y=z>>3,w=u.ra[Y],D&&(v=z,V=u,V.L!=v>>6&&(V.L=v>>6,H=m(V,274),V.PQ=K0(15,255,V.Y,V.L,[0,0,H[1],H[2]])),w^=u.PQ[Y&E]),q|=(w>>8-(R|0)-(x|0)&(1<<x)-1)<<(J|0)-(x|0),J-=x,z+=x;return(n=q,y)(u,(Z|0)+(Q|0),490),n},En=typeof Object.defineProperties=="function"?Object.defineProperty:function(u,Q,D,Y){{Y=37;while(Y!=32)if(Y==37)Y=u==Array.prototype||u==Object.prototype?36:8;else{if(Y==8)return u[Q]=D.value,u;if(Y==36)return u}}},K0=function(u,Q,D,Y,w,v,J,n){for(J=w[3]|(n=w[2]|(v=0,0),0);v<u;v++)Y=Y>>>8|Y<<24,Y+=D|0,J=J>>>8|J<<24,D=D<<3|D>>>29,Y^=n+2167,J+=n|0,D^=Y,J^=v+2167,n=n<<3|n>>>29,n^=J;return[D>>>24&Q,D>>>16&Q,D>>>8&Q,D>>>0&Q,Y>>>24&Q,Y>>>16&Q,Y>>>8&Q,Y>>>0&Q]},IZ=function(u,Q,D,Y,w,v,J,n,H,z){for(u.Bm=m6(41,u.A,(u.zJ=(u.EI=Tu,eF),u.lw=u[Sz],{get:function(){return this.concat()}})),u.Yh=hl[u.A](u.Bm,{value:{value:{}}}),n=[],H=0;H<294;H++)n[H]=String.fromCharCode(H);u.n8=false,(u.jl=0,u).J=(u.t0=25,u.N=(u.bO=void 0,false),u.da=0,u.EW=(u.yP=false,[]),false);while(0==![undefined])if(u.T=u,[])break;if((u.oh=(u.Ac=(u.H=0,(u.I=void 0,u.G=0,u.o=null,u.uO=(u.iO=void 0,0),u).QP=(z=(u.aM=J,window.performance||{}),(u.hc=!(u.p7=[],u.WQ=0,u.kB=(u.PQ=void 0,0),((u.ra=(u.cm=D,[]),u.mM=[],u).ej=(u.Y=void 0,u.h0=0,u.TJ=8001,function(b){return s4.call(this,33,8,b)}),u).K=1,1),u.xB=false,u.C=[],(u.s=void 0,u.L=void 0,u).h=void 0,u).OW=[],[]),z.timeOrigin||(z.timing||{}).navigationStart||0),u.W=[],0),Y&&Y.length==2)&&(u.p7=Y[1],u.mM=Y[0]),Q)try{u.iO=JSON.parse(Q)}catch(b){u.iO={}}if(![]==(ZY(0,(l(280,u,(u.Qg=(l(133,u,66,(l(325,(l(459,(l(29,u,66,(l(46,u,(l(138,u,70,(L(373,u,(l(106,u,((l(502,(l(123,u,(l(224,(l(226,(l(408,u,(l((L(68,(L(114,(l(427,u,(l(340,u,75,(l(180,u,67,(y(u,(l(292,u,(B((y(u,(l(309,u,64,(L(76,u,(l(310,(l(28,u,(l((l(497,u,77,(l(57,u,(l(265,(l(281,(L(302,u,(L(268,(B((L(18,u,(B(492,((B(156,0,(y(u,(l(82,(y(u,0,(l(193,u,(B((y(u,(l(51,u,73,(l(482,u,(l(475,u,65,function(b,x,V,Z,R,E,q,h,r){{r=64;while(r!=89)r==40?r=R--?65:7:r==68?r=40:r==30?r=40:r==65?(E=(Z=Ks(true,38,b,128),-~(E&Z)+-2-~(E|Z))%q,x.push(h[E]),r=68):r==7?(B(V,x,b),r=89):r==64&&(V=F(b,8),R=Ks(true,33,b,128),x=[],h=I(b,159),E=0,q=h.length,r=30)}}),77),function(b,x,V,Z,R,E,q,h,r,A){for(A=27;A!=46;)A==11?(Z++,A=36):A==3?A=36:A==2?(R+=String.fromCharCode((r=E[Z],-121+(r|121)+(~r&121))),A=11):A==40?(L(x,b,h[R]),A=46):A==36?A=Z<E.length?2:40:A==27&&(q=W(5,b),V=F(b,7),x=W(5,b),h=m(b,q),E=k(V,b),R="",Z=0,A=3)}),function(b,x,V,Z,R,E,q,h,r,A){for(A=1;A!=57;)A==1?(r=W(17,b),h=W(13,b),x=W(55,b),V=k(r,b),E=k(h,b),q="",R=0,A=48):A==72?(y(b,q in E|0,x),A=57):A==87?(R++,A=93):A==93?A=R<V.length?74:72:A==74?(q+=String.fromCharCode((Z=V[R],-1+(~Z&121)-(~Z|121))),A=87):A==48&&(A=93)})),0),490),72),0,u),u.iw=0,78),function(b){Ks(true,16,4,2,b)}),185)),u),71,function(b){WG(b,1)}),aZ(4)),230),u)),l)(214,u,68,function(b,x,V){(x=k((V=F(b,7),V),b.T),x)[0].removeEventListener(x[1],x[2],cK)}),e),u),[])),250),[0,0,0],u),u),[2048]),[])),u),64,function(b){BG(b,3)}),u),67,function(b,x,V,Z,R,E,q,h,r,A,X,U,d,c,a){for(a=59;a!=83;)if(a==82)a=X<r?51:83;else if(a==51)Z(A.slice(X,(X|0)+(c|0)),R),a=57;else if(a==2)a=82;else if(a==57)X+=c,a=82;else if(a==20){for(E in d=[],A)d.push(E);a=(A=d,61)}else a==81?(h=F(b,5),q=W(45,b),U=W(47,b),V=F(b,3),A=k(h,b),R=I(b,V),c=m(b,U),Z=I(b,q),a=68):a==68?a=XB("array",A,"object")=="object"?20:61:a==36?(c=c>0?c:1,r=A.length,X=0,a=2):a==61?a=b.T==b?36:83:a==59&&(a=m6(90,true,2,true,x,b)?83:81)}),69),function(b,x){XM(268,104,(x=I(b,W(45,b)),b.T),0,490,x)}),y(u,[],254),function(b,x,V,Z,R,E,q,h,r,A){for(A=38;A!=78;)A==38?A=m6(88,false,2,true,x,b)?78:83:A==83&&(h=$L(13,3,b.T,1),V=h.X2,r=h.jj,q=h.UW,Z=h.i,E=Z.length,R=E==0?new r[q]:E==1?new r[q](Z[0]):E==2?new r[q](Z[0],Z[1]):E==3?new r[q](Z[0],Z[1],Z[2]):E==4?new r[q](Z[0],Z[1],Z[2],Z[3]):2(),L(V,b,R),A=78)})),236),u,72,function(b,x,V,Z,R,E,q,h,r){for(r=79;r!=30;)r==93?r=q--?16:88:r==79?(Z=W(37,b),q=Ks(true,37,b,128),E="",V=m(b,159),x=V.length,h=0,r=94):r==16?(h=(R=Ks(true,35,b,128),2*(h&R)+(h&~R)+(~h&R))%x,E+=n[V[h]],r=6):r==94?r=93:r==88?(L(Z,b,E),r=30):r==6&&(r=93)}),66),function(b,x,V,Z){x=$f(true,(Z=W(5,b),b),8),V=F(b,7),L(V,b,I(b,Z)>>>x)}),u),79,function(b,x,V,Z,R,E){y((x=m(b,(Z=I(b,(V=W(33,(R=F(b,6),b)),E=W(15,b),R)),V)),b),Z in x|0,E)}),aZ(4))),function(b,x,V){(V=W(15,(x=F(b,3),b)),L)(V,b,""+m(b,x))})),[]),314),267),u,u),75),function(b,x,V,Z,R){y(b,(x=I(b,(R=I((Z=F(b,(V=F(b,7),3)),b),V),Z)),x+R),Z)}),{}),244),function(b,x){(x=W(49,b),L)(x,b,[])})),u.Jc=0,function(b,x,V,Z,R){{R=85;while(R!=94)R==92?(V=W(13,b),Z=F(b,3),L(Z,b,function(E){return eval(E)}(FM(I(b.T,V)))),R=94):R==85&&(R=m6(91,false,2,true,x,b)?94:92)}})),65),function(b){BG(b,4)}),u),604),u),aZ(4)),464),u,73,function(){}),79),function(b,x,V,Z,R,E,q,h,r,A,X){{X=96;while(X!=94)X==99?(q=W(6,2,false,b,r,Z,1,E,R),E.addEventListener(R,q,cK),k(302,b).push(function(){E.removeEventListener(R,q,cK)}),L(156,b,[E,R,q]),X=94):X==96?(A=W(13,b),h=W(49,b),V=F(b,5),x=W(17,b),r=m(b,V),R=I(b,h),E=k(A,b.T),Z=m(b,x),X=55):X==55&&(X=E!==0?99:94)}}),u),71,function(b){WG(b,4)}),u),70,function(b,x,V,Z,R,E){{E=9;while(E!=32)E==21?E=b.T==b||V==b.ej&&Z==b?27:32:E==27?(L(R.X2,b,V.apply(Z,R.i)),b.jl=b.X(),E=32):E==37?(R=$L(13,3,b,1),V=R.UW,Z=R.jj,E=21):E==9&&(E=m6(89,false,2,true,x,b)?32:37)}}),74),function(b,x,V,Z,R,E){V=I(b,(E=m(b,(R=W(23,(Z=(x=W(37,b),W)(5,b),b)),Z)),x))==E,L(R,b,+V)}),u),78,function(b,x,V,Z,R,E){{E=25;while(E!=39)E==50?(R++,E=46):E==25?(x=W(5,b),V=Ks(true,34,b,128),Z=[],R=0,E=93):E==46?E=R<V?35:53:E==93?E=46:E==35?(Z.push($f(true,b,8)),E=50):E==53&&(B(x,Z,b),E=39)}}),B)(40,[],u),74),function(b,x,V,Z,R,E,q,h){if(q=W(55,b),2)Z=F(b,5);y(b,W(8,2,(R=m(b,(V=m(b,(E=(x=(h=F(b,8),W)(47,b),I)(b,x),h)),Z)),false),b,R,V,E),q)}),[165,0,0])),function(b,x,V,Z,R,E,q,h,r,A,X,U,d,c,a,p,G$,vK,K){for(K=46;K!=16;)K==80?K=12:K==2?(Z=vK(1),A.push(Z),R+=Z?0:1,K=95):K==46?(vK=function(S,O){for(;V<S;)h|=$f(true,b,8)<<V,V+=8;return h>>=(O=h&((V-=S,1)<<S)-1,S),O},U=F(b,6),V=h=0,G$=(x=vK(3),2*(x&1)-1-(~x^1)),c=vK(5),A=[],r=R=0,K=90):K==91?K=d<c?72:84:K==10?K=12:K==55?(A[q]&&(p[q]=W(45,b)),K=65):K==90?K=6:K==6?K=r<c?2:63:K==28?(l(U,b,64,function(S,O,HK,ME,R_,N){for(N=8;N!=49;)N==60?N=O>=HK.length?97:44:N==8?(R_=0,HK=[],ME=[],N=14):N==21?(O=p[R_],N=7):N==70?(S.s=F(S,10,a.slice()),S.I=F(S,9,ME),N=49):N==14?N=2:N==78?(ME.push(O),N=66):N==7?N=A[R_]?78:75:N==2?N=R_<c?21:70:N==66?(R_++,N=2):N==35?N=60:N==44?(O=HK[O],N=78):N==75?N=60:N==97&&(HK.push(F(S,6)),N=35)}),K=16):K==1?K=q<c?55:34:K==65?(q++,K=1):K==95?(r++,K=6):K==34?(X=G$,a=[],K=10):K==72?(A[d]||(p[d]=vK(E)),K=68):K==96?K=91:K==68?(d++,K=91):K==84?(q=0,K=40):K==43?(a.push(m(b,W(55,b))),K=80):K==40?K=1:K==63?(E=((R|0)-1).toString(2).length,p=[],d=0,K=96):K==12&&(K=X--?43:28)})),65),function(b,x,V,Z,R){(Z=(x=m(b,(V=W(55,(R=W(17,b),b)),R))!=0,k(V,b)),x)&&L(490,b,Z)}),function(b,x,V,Z){L((Z=(x=(V=W(47,b),W(15,b)),W(15,b)),Z),b,k(V,b)||m(b,x))})),(new AM("Submit")).dispose(),u),68,function(b,x,V,Z,R,E){V=I(b,(Z=I(b,(x=F(b,(E=W(45,b),8)),R=W(49,b),E)),x)),L(R,b,Z[V])}),u),69,function(b,x,V,Z,R,E,q,h){{h=18;while(h!=94)h==18?(R=W(37,b),Z=W(23,b),q=W(47,b),h=50):h==50?h=b.T==b?0:94:h==65?(b.L=void 0,h=30):h==30?h=E==2?11:94:h==0?(E=I(b,Z),V=m(b,R),x=m(b,q),V[E]=x,h=63):h==11?(b.Y=M(b,32,false),b.L=void 0,h=94):h==63&&(h=R==274?65:94)}}),function(b,x,V,Z,R){for(R=59;R!=52;)R==3?R=Z?49:75:R==75?(B(490,b.G,b),R=52):R==15?R=2:R==77?(Z[18]=b.C[18],Z[268]=b.C[268],b.C=Z,R=52):R==49?(x=$f(true,b,8),R=15):R==72?(x--,R=2):R==2?R=x>0?18:77:R==18?(V=W(33,b),Z[V]=b.C[V],R=72):R==59&&(Z=b.QP.pop(),R=3)})),0),72),function(b,x,V,Z,R){y((R=XB("array",(Z=I(b,(V=F(b,(x=W(33,b),6)),x)),Z),"object"),b),R,V)}),22),u,[il]),0))ZY(0,14,u,[ia,w]);G(16,254,(ZY(0,23,u,[kL,v]),true),true,u)},u3=function(u,Q,D,Y,w){return jz.call(this,8,48,u,Q,D,Y,w)},BG=function(u,Q,D,Y,w,v,J){(D=m(u,(v=(Y=(J=(Q|(w=Q&4,0))-~(Q&3)+~(Q|3)+(~Q&3),F(u,3)),F(u,5)),Y)),w&&(D=f0(224,""+D)),J&&y9(2,P(2,D.length),v,u),y9)(2,D,v,u)},qE=function(u,Q){while([]){return ZY.call(this,u,3,Q);if("E")break}},L0=function(){return Ls.call(this,2,48)},t,$f=function(u,Q,D){return Q.s?FB(Q,Q.I):M(Q,D,u)},n0=function(){return bl.call(this,14,3)},la=function(u,Q,D,Y,w,v,J,n){if(!D.h){D.WQ++;try{for(w=(J=(v=void 0,0),D).G;--Q;)try{if(n=void 0,D.s)v=FB(D,D.s);else{if((J=m(D,490),J)>=w)break;v=k((n=F(D,(y(D,J,72),6)),n),D)}v&&v[C0]&2048?v(D,Q):Gu(0,[gX,21,n],D,Y),m6(92,false,2,false,Q,D)}catch(H){m(D,u)?Gu(22,H,D,Y):y(D,H,u)}while(!Q){switch(!D.n7){case 0==![""]:void(!(!""!=!false)==!"").true;break;case true==[]:la(114,729113759829,(D.WQ--,D),268);return;break}if(!""==(Gu(0,[gX,33],D,Y),!false))break}}catch(H){try{Gu(22,H,D,Y)}catch(z){G(41,0,z,D)}}D.WQ--}},b3=function(u,Q,D,Y,w,v,J,n,H,z,b,x){{b=98;while(b!=19)if(b==2)z++,b=30;else if(b==91){a:{if(n&&typeof n.length=="number"){if(BK(58,31,"object",n)){H=typeof n.item=="function"||typeof n.item==Q;break a}if(typeof n==="function"){H=typeof n.item=="function";break a}}H=false}Yf(75,48,u,v,x,H?m6(16,n,u):n),b=2}else b==98?(x=function(V){V&&w.appendChild(typeof V==="string"?J.createTextNode(V):V)},z=1,b=71):b==30?b=z<Y.length?72:19:b==73?b=!fs(50,"object",6,D,"number",n)||BK(58,34,"object",n)&&n.nodeType>u?49:91:b==71?b=30:b==72?(n=Y[z],b=73):b==49&&(x(n),b=2)}},jF=function(u,Q,D,Y,w,v){return U4.call(this,w,Q,v,31,D,u,Y)},wG=function(u,Q,D,Y){try{Y=u[(-~(Q&2)+-2-~Q+(~Q&2))%3],u[Q]=(u[Q]|0)-(u[(-2-3*~(Q|1)-(~Q&1)+2*(~Q|1))%3]|0)-(Y|0)^(Q==1?Y<<D:Y>>>D)}catch(w){throw w;}},zu=function(){return G.call(this,48)},XM=function(u,Q,D,Y,w,v){while(5)if(D.QP.length>Q?Gu(Y,[gX,36],D,u):(D.QP.push(D.C.slice()),D.C[w]=void 0,L(w,D,v)),true)break},B=function(u,Q,D){switch(!(u==490||u==72)){case ![]==(true==![]):while(D.n8&&u!=274){return;if({})break}u==373||u==76||u==314||u==230||u==18||u==40||u==254||u==250||u==68||u==268?D.C[u]||(D.C[u]=Q9(D,Q,6,17,30,u)):D.C[u]=Q9(D,Q,6,18,41,u);break;case false:D.C[u]?D.C[u].concat(Q):D.C[u]=F(D,12,Q);break}u==274&&(D.Y=M(D,32,false),D.L=void 0)},Qu=function(){return xf.call(this,17,7)},g=function(u,Q,D,Y,w,v,J){J=this;try{IZ(this,w,v,Y,Q,D,u)}catch(n){G(27,0,n,this),D(function(H){H(J.h)})}},D5=function(u){return kf.call(this,3,3,u)},oZ=m6(12,"Math",0,"object",this),e=(VR(8,".",null,1,0,"Symbol",function(u,Q,D,Y,w,v){for(w=70;w!=67;){if(w==23)return u;if(w==92)return v.prototype.toString=function(){return this.uw},D="jscomp_symbol_"+(Math.random()*1E9>>>0)+"_",Q=0,Y;w==85?w=u?23:92:w==70&&(v=function(J,n){En((this.uw=J,this),"description",{configurable:true,writable:true,value:n})},Y=function(J,n){for(n=77;n!=36;){if(n==46)return new v(D+(J||"")+"_"+Q++,J);if(n==84)throw new TypeError("Symbol is not a constructor");n==77&&(n=this instanceof Y?84:46)}},w=85)}}),this||self),WK="closure_uid_"+(Math.random()*1E9>>>0),NE=0,V9,YL=function(u,Q,D,Y,w,v){for(Y=91,v=78;;)try{if(Y==29)break;else if(Y==43)D=false,u=Object.defineProperty({},"passive",{get:function(){D=true}}),Y=38;else if(Y==91)Y=e.addEventListener&&Object.defineProperty?43:66;else if(Y==55)v=78,Y=53;else{if(Y==53)return v=78,D;if(Y==38)v=7,Q=function(){},e.addEventListener("test",Q,u),e.removeEventListener("test",Q,u),Y=53;else if(Y==66)return false}}catch(J){if(v==78)throw J;v==7&&(w=J,Y=55)}}(),ps="closure_listenable_"+(((Cs(22,28,2,rZ,(a_.prototype.Z=function(u){for(u=19;u!=74;)u==41?(this.ga.shift()(),u=4):u==85?u=this.ga.length?41:74:u==4?u=85:u==36?u=85:u==19&&(u=this.ga?36:74)},a_.prototype[(qE.prototype.preventDefault=function(){this.defaultPrevented=true},qE).prototype.stopPropagation=function(){this.Te=true},(a_.prototype.dispose=function(u){{u=50;while(u!=31)u==80?(this.P=true,this.Z(),u=31):u==50&&(u=this.P?31:80)}},a_.prototype).P=false,Symbol.dispose]=function(){this.dispose()},qE)),rZ.prototype.stopPropagation=function(){rZ.j.stopPropagation.call(this),this.U.stopPropagation?this.U.stopPropagation():this.U.cancelBubble=true},rZ).prototype.preventDefault=function(u){u=(rZ.j.preventDefault.call(this),this.U),u.preventDefault?u.preventDefault():u.returnValue=false},Math.random()*1E6)|0),PG="constructor hasOwnProperty isPrototypeOf propertyIsEnumerable toLocaleString toString valueOf".split(" "),Zi=0,PK="closure_lm_"+((yR.prototype.add=((yR.prototype.HQ=function(u,Q,D,Y,w,v){return((v=this.B[u.toString()],w=-1,v)&&(w=jz(8,5,0,Q,v,D,Y)),w>-1)?v[w]:null},yR.prototype).remove=function(u,Q,D,Y,w,v,J,n){{n=8;while(n!=45){if(n==32)return false;if(n==50)delete this.B[w],this.XH--,n=63;else if(n==15)n=J>-1?64:32;else if(n==4)v=this.B[w],J=jz(8,3,0,Q,v,D,Y),n=15;else{if(n==63)return true;if(n==64)ul(true,7,v[J]),Array.prototype.splice.call(v,J,1),n=77;else if(n==8)w=u.toString(),n=75;else{if(n==11)return false;n==77?n=v.length==0?50:63:n==75&&(n=w in this.B?4:11)}}}}},function(u,Q,D,Y,w,v,J,n,H,z){{z=7;while(z!=73)if(z==83)n=new Mm(w,Q,this.src,v,!!Y),n.sW=D,H.push(n),z=16;else{if(z==16)return n;z==7?(v=u.toString(),H=this.B[v],z=15):z==74?(J=jz(8,6,0,Q,H,Y,w),z=45):z==45?z=J>-1?51:83:z==41?z=D?16:87:z==51?(n=H[J],z=41):z==87?(n.sW=false,z=16):z==15?z=H?74:24:z==24&&(H=this.B[v]=[],this.XH++,z=74)}}}),yR.prototype).hasListener=function(u,Q,D,Y,w){return DY(37,false,(w=(Y=u!==(D=Q!==void 0,void 0))?u.toString():"",true),16,this.B,function(v,J,n){{n=38;while(n!=48){if(n==76)return true;if(n==38)J=0,n=35;else{if(n==13)return false;n==21?n=Y&&v[J].type!=w||D&&v[J].capture!=Q?59:76:n==35?n=0:n==0?n=J<v.length?21:13:n==59&&(++J,n=0)}}}})},Math.random()*1E6|0),o_={},wX=0,tl="__closure_events_fn_"+(Math.random()*1E9>>>0);if((t=((Cs(22,16,2,n0,a_),n0).prototype[ps]=true,n0.prototype),t.VP=function(u){this.A0=u},t).addEventListener=function(u,Q,D,Y){s4(33,18,"object",false,Y,Q,u,this,D)},t.removeEventListener=function(u,Q,D,Y){O4(0,14,"object",Q,Y,D,u,this)},[])t.dispatchEvent=function(u,Q,D,Y,w,v,J,n,H,z,b,x){{x=43;while(x!=25)if(x==51)x=z.Te?18:92;else if(x==99)x=81;else if(x==84)x=typeof z==="string"?24:62;else if(x==33)w--,x=57;else if(x==43)n=this.A0,x=71;else if(x==39)x=59;else if(x==15)z=u,b=this.L7,H=z.type||z,Y=Q,x=84;else if(x==24)z=new qE(z,b),x=60;else if(x==78)x=57;else if(x==71)x=n?68:15;else if(x==26)z.target=z.target||b,x=60;else if(x==53)D=z,z=new qE(H,b),sn(z,D),x=60;else if(x==60)J=true,x=48;else if(x==97)v=z.currentTarget=Y[w],J=RZ(5,true,z,v,H,false)&&J,x=7;else if(x==9)v=z.currentTarget=Y[w],J=RZ(6,true,z,v,H,true)&&J,x=33;else if(x==81)x=!z.Te&&w<Y.length?97:74;else if(x==18)x=Y?20:74;else if(x==48)x=Y?63:51;else if(x==94)Q.push(n),x=3;else if(x==7)w++,x=81;else if(x==3)n=n.A0,x=59;else if(x==59)x=n?94:15;else if(x==92)v=z.currentTarget=b,J=RZ(8,true,z,v,H,true)&&J,z.Te||(J=RZ(7,true,z,v,H,false)&&J),x=18;else if(x==62)x=z instanceof qE?26:53;else if(x==20)w=0,x=99;else if(x==57)x=!z.Te&&w>=0?9:51;else{if(x==74)return J;x==68?(Q=[],x=39):x==63&&(w=Y.length-1,x=78)}}};t.Z=(t.hasListener=function(u,Q){return this.u.hasListener(u!==void 0?String(u):void 0,Q)},t.HQ=function(u,Q,D,Y){return this.u.HQ(String(u),Q,D,Y)},function(){n0.j.Z.call(this),this.u&&E4(94,true,0,17,this.u),this.A0=null});var JM;(((((t=("ARTICLE SECTION NAV ASIDE H1 H2 H3 H4 H5 H6 HEADER FOOTER ADDRESS P HR PRE BLOCKQUOTE OL UL LH LI DL DT DD FIGURE FIGCAPTION MAIN DIV EM STRONG SMALL S CITE Q DFN ABBR RUBY RB RT RTC RP DATA TIME CODE VAR SAMP KBD SUB SUP I B U MARK BDI BDO SPAN BR WBR NOBR INS DEL PICTURE PARAM TRACK MAP TABLE CAPTION COLGROUP COL TBODY THEAD TFOOT TR TD TH SELECT DATALIST OPTGROUP OPTION OUTPUT PROGRESS METER FIELDSET LEGEND DETAILS SUMMARY MENU DIALOG SLOT CANVAS FONT CENTER ACRONYM BASEFONT BIG DIR HGROUP STRIKE TT".split(" ").concat(["BUTTON","INPUT"]),zu.prototype),t.F=function(u){return typeof u==="string"?this.el.getElementById(u):u},t.getElementsByTagName=function(u,Q){return(Q||this.el).getElementsByTagName(String(u))},t.createElement=function(u,Q,D){return((Q=String((D=this.el,u)),D).contentType==="application/xhtml+xml"&&(Q=Q.toLowerCase()),D).createElement(Q)},t).createTextNode=function(u){return this.el.createTextNode(String(u))},t).appendChild=function(u,Q){u.appendChild(Q)},t.append=function(u,Q){b3(0,"string","array",arguments,u,"",u.nodeType==9?u:u.ownerDocument||u.document)},t).canHaveChildren=function(u,Q){for(Q=28;Q!=8;){if(Q==86)return false;if(Q==28)Q=u.nodeType!=1?86:57;else if(Q==57){switch(u.tagName){case "APPLET":case "AREA":case "BASE":case "BR":case "COL":case "COMMAND":case "EMBED":case "FRAME":case "HR":case "IMG":case "INPUT":case "IFRAME":case "ISINDEX":case "KEYGEN":case "LINK":case "NOFRAMES":case "NOSCRIPT":case "META":case "OBJECT":case "PARAM":case "SCRIPT":case "SOURCE":case "STYLE":case "TRACK":case "WBR":return false}return true}}},t.removeNode=D5,t).contains=function(u,Q,D){{D=98;while(D!=57)if(D==98)D=u&&Q?99:31;else{if(D==78)return u==Q||!!(u.compareDocumentPosition(Q)&16);if(D==80)D=40;else if(D==86)Q=Q.parentNode,D=80;else if(D==26)D=40;else{if(D==81)return Q==u;if(D==51)return u==Q||u.contains(Q);if(D==99)D=u.contains&&Q.nodeType==1?51:7;else{if(D==31)return false;D==7?D=typeof u.compareDocumentPosition!="undefined"?78:26:D==40&&(D=Q&&u!=Q?86:81)}}}}},ul(rX,78),rX.prototype).gp="";while(2)if(rX.prototype.yg=0,{})break;(((t=(Cs(22,12,2,ns,n0),ns).prototype,t.Wm=rX.p8(),t).F=function(){return this.v},t.getParent=function(){return this.qk},t.Z=function(u){{u=79;while(u!=78)u==80?u=this.C8?19:3:u==19?(this.C8.dispose(),delete this.C8,u=3):u==79?(this.vQ&&this.D(),u=80):u==3&&(fs(50,this,22,function(Q){Q.dispose()}),!this.MI&&this.v&&D5(this.v),this.qk=this.Zt=this.v=this.Sl=null,ns.j.Z.call(this),u=78)}},t.VP=function(u,Q){for(Q=15;Q!=80;){if(Q==23)throw Error("Method not supported");Q==50?(ns.j.VP.call(this,u),Q=80):Q==15&&(Q=this.qk&&this.qk!=u?23:50)}},t).D=function(){(fs(50,this,23,function(u){u.vQ&&u.D()}),this.C8&&E4(94,true,0,18,this.C8),this).vQ=false},t).removeChild=function(u,Q,D,Y,w,v,J,n,H,z,b,x,V){{V=36;while(V!=25)if(V==51)n=u,V=0;else if(V==5)w=x,V=95;else if(V==58)V=u?39:99;else{if(V==99)throw Error("Child is not in parent component");if(V==82)D=this.Sl,v=(D!==null&&w in D?D[w]:void 0)||null,V=59;else if(V==56)H=u,b=u.Wm,Y=b.gp+":"+(b.yg++).toString(36),J=H.rp=Y,V=97;else if(V==63)V=Q?32:51;else if(V==26)V=w&&u?38:58;else if(V==1)v=null,V=59;else{if(V==52)throw Error("Unable to set parent component");if(V==0)V=n==null?52:41;else if(V==95)V=this.Sl&&w?82:1;else if(V==40)V=(J=u.rp)?97:56;else if(V==41)n.qk=null,ns.j.VP.call(n,null),V=58;else if(V==97)x=J,V=5;else{if(V==39)return u;V==84?(x=u,V=5):V==38?(z=this.Sl,w in z&&delete z[w],VR(18,0,u,this.Zt),V=63):V==59?(u=v,V=26):V==36?V=u?72:58:V==72?V=typeof u==="string"?84:40:V==32&&(u.D(),u.v&&D5(u.v),V=51)}}}}};var YF,jb={button:"pressed",checkbox:"checked",menuitem:"selected",menuitemcheckbox:"checked",menuitemradio:(t=(ul(Qu,70),Qu.prototype),t.Mk=function(u){return u.F()},"checked"),radio:"checked",tab:"selected",treeitem:"selected"},Jl=(ul(L0,(Cs(22,16,2,(t.IM=((t.mH=function(u,Q,D,Y){(Y=u.F?u.F():u)&&(D?u3:qm)(Y,[Q])},t).FH=(t.g=function(u,Q,D,Y,w,v,J){for(J=14;J!=49;)J==67?J=this.K8?80:36:J==14?(v=Q.F(),J=99):J==36?(w=this.Dt(),w.replace(/\\xa0|\\s/g," "),this.K8={1:w+"-disabled",2:w+"-hover",4:w+"-active",8:w+"-selected",16:w+"-checked",32:w+"-focused",64:w+"-open"},J=80):J==80?((Y=this.K8[u])&&this.mH(Q,Y,D),this.IM(v,u,D),J=49):J==99&&(J=v?67:49)},function(u,Q,D,Y,w,v,J,n,H){for(J=(n=77,20);;)try{if(n==50)break;else n==17?(D.tabIndex=0,n=50):n==61?(D.tabIndex=-1,D.removeAttribute("tabIndex"),n=50):n==55?(J=20,n=66):n==49?(u.f8&4&&I_(u,17,4,1)&&u.setActive(false),u.f8&32&&I_(u,48,32,1)&&RZ(24,32,u,32,false)&&u.g(false,32),n=48):n==48?n=(w=v.hasAttribute("tabindex"))?85:80:n==28?(D=v,n=69):n==12?(J=20,n=55):n==66?n=u.S&32?49:48:n==85?(Y=v.tabIndex,w=typeof Y==="number"&&Y>=0&&Y<32768,n=80):n==88?n=!Q&&u.S&32?46:48:n==69?n=Q?17:61:n==46?(J=27,v.blur(),n=55):n==80?n=w!=Q?28:50:n==77&&(n=I_(u,49,32,1)&&(v=u.Mk())?88:50)}catch(z){if(J==20)throw z;J==27&&(H=z,n=12)}}),function(u,Q,D,Y,w,v,J,n){(w=(Y=(YF||(YF={1:"disabled",8:"selected",16:"checked",64:"expanded"}),YF[Q]),u.getAttribute("role")||null))?(J=jb[w]||Y,v=Y=="checked"||Y=="selected"?J:Y):v=Y;while(NaN!==Number(undefined))if((n=v)&&dZ("hidden",u,"none",9," ",D,n),![]!=true)break}),t.Dt=function(){return"goog-control"},L0),Qu),71)),{});(((((((t=(Cs((L0.prototype.Dt=(L0.prototype.IM=function(u,Q,D){switch(Q){case 8:case 16:dZ("hidden",u,"none",3," ",D,"pressed");break;default:case 64:case 1:L0.j.IM.call(this,u,Q,D)}},function(){while(0==![]){return"goog-button";if([])break}}),22),28,2,vG,ns),vG).prototype,t.mH=function(u,Q,D){for(D=75;D!=98;)D==10?(this.m=null,D=6):D==82?D=u&&this.m&&VR(26,0,u,this.m)?0:98:D==75?D=Q?54:82:D==0?D=this.m.length==0?10:6:D==54?D=u?93:98:D==6?(this.l.mH(this,u,false),D=98):D==93&&(this.m?kf(3,11,0,this.m,u)>=0||this.m.push(u):this.m=[u],this.l.mH(this,u,true),D=98)},t.bw=0,t.S=0,t.D=function(){((vG.j.D.call(this),this.YB)&&this.YB.detach(),this.isVisible()&&this.isEnabled())&&this.l.FH(this,false)},t).GJ=true,t).Z=function(u){for(u=65;u!=18;)u==17?(this.YB.dispose(),delete this.YB,u=1):u==65?(vG.j.Z.call(this),u=47):u==1?(delete this.l,this.m=null,u=18):u==47&&(u=this.YB?17:1)},t.f8=255,t).m=null,t.Mk=function(){return this.l.Mk(this)},t.Ih=39,t).isVisible=function(){return this.GJ},t).isEnabled=function(){while(true){return!(this.S&1);if(!null)break}},t.isActive=function(){return!!(this.S&4)},t.setActive=function(u){RZ(25,32,this,4,u)&&this.g(u,4)},t).getState=function(){return this.S},t).g=function(u,Q,D,Y,w,v,J){for(J=44;J!=8;)J==19?(this.isVisible()&&this.l.FH(this,Y),this.g(!Y,1,true),J=8):J==12?J=Y?19:61:J==53?(this.l.g(Q,this,u),this.S=u?this.S|Q:(w=this.S,~Q- -1+(w|~~Q)),J=8):J==44?J=D||Q!=1?66:75:J==75?(Y=!u,v=this.getParent(),J=59):J==59?J=v&&typeof v.isEnabled=="function"&&!v.isEnabled()||!RZ(26,32,this,1,!Y)?8:12:J==66?J=I_(this,33,Q,1)&&u!=!!(this.S&Q)?53:8:J==61&&(this.setActive(false),RZ(27,32,this,2,false)&&this.g(false,2),J=19)};for(true;typeof vG!=="function";![]==0){throw Error("Invalid component class "+vG);if(![(!false==!"").true]==Number())break}for(false;typeof Qu!=="function";undefined){throw Error("Invalid renderer class "+Qu);if(true)break}var vp=xf(17,16,vG),cK={passive:true,capture:(E4(94,function(){return new AM(null)},"goog-button",((Cs(22,12,2,(((ul(xL,(Cs(22,(E4((Jl[vp]=Qu,94),function(){return new vG(null)},"goog-control",5),32),2,xL,L0),77)),xL).prototype.IM=function(){},xL).prototype.FH=function(){},xL.prototype.g=function(u,Q,D,Y,w){for(w=15;w!=77;)w==78?w=Y&&u==1?40:77:w==40?(Y.disabled=D,w=77):w==15&&(xL.j.g.call(this,u,Q,D),Y=Q.F(),w=78)},AM),vG),AM).prototype.Z=function(){delete (AM.j.Z.call(this),this).tc,delete this.ah},9)),true)},Al=e.requestIdleCallback?function(u){requestIdleCallback(function(){u()},{timeout:4})}:e.setImmediate?function(u){setImmediate(u)}:function(u){setTimeout(u,0)},mN=String.fromCharCode(105,110,116,101,103,67,104,101,99,107,66,121,112,97,115,115),T$=[],kL=[],il=[],ia=[];g.prototype.oM="toString";while(0==![undefined])if(g.prototype.NI=void 0,[])break;var gX=(g.prototype.xh=void 0,{}),gZ=(g.prototype.n7=false,[]),Sz=[],ll=[],C0=[];while(0===-0)if(![]==(tM,false==null))break;var hl=(((((aZ,function(){})(wG),function(){})(hM),function(){})(Un),function(){})(dX),g.prototype.A="create",gX.constructor),ua=(((t=g.prototype,t).J0=function(u,Q,D,Y,w,v){return W.call(this,66,u,Q,D,Y,w,v)},t.Vg=0,t).kh=function(){return bl.call(this,14,16)},void 0);if(0===-((t.X=(window.performance||{}).now?function(){return this.Ac+window.performance.now()}:function(){return+new Date},t).Rh=function(){return Ls.call(this,2,26)},Number()))t.OI=function(u,Q,D,Y,w,v){return HG.call(this,24,18,u,Q,D,Y,w,v)};(((t=(t.Hm=function(u,Q,D,Y){return I_.call(this,Q,3,D,u,Y)},t.F2=function(u,Q,D,Y,w,v,J,n,H,z){while(0===-0){return I_.call(this,Q,28,D,u,Y,w,v,J,n,H,z);if(15)break}},g).prototype,t).R=function(u,Q){return ua=function(){return Q==u?73:53},u=(Q={},{}),function(D,Y,w,v,J,n,H,z,b,x,V,Z,R,E,q,h,r,A,X,U,d,c,a,p,G$,vK,K,S,O,HK,ME,R_,N,Di,f,Jj,wZ,cG,T,nD){wZ=(f=(T=41,8),undefined);{Jj=false;while(![]==0)try{if(f==80)break;else if(f==32)f=R==ia?46:91;else if(f==22)f=w.length>4?59:49;else if(f==66)h=Z.value,f=30;else if(f==20)f=R==gZ?86:82;else if(f==51)C(373,this,P(2,w.length).concat(w),153),f=49;else if(f==26)f=Z.done?83:66;else if(f==87)f=98;else if(f==77)T=40,a=aZ(2).concat(I(this,373)),a[1]=(r=a[0],-(r&3)-~(r&3)+-2-(~r^3)),a[3]=(A=a[1],v=G$[0],-1+(A&~v)-(A|~v)),a[4]=a[1]^G$[1],J=this.Sj(a),f=23;else if(f==38)T=40,la(114,8001,this,268),f=15;else if(f==23)f=J?88:13;else if(f==24)wZ!==undefined?(f=wZ,wZ=undefined):f=80;else{if(f==90)return Di;if(f==7)T=40,R=D[0],f=32;else if(f==52)f=b<a.length?19:53;else if(f==67)f=R==C0?65:15;else if(f==45)w=w.slice(0,1E6),C(373,this,[],250),C(373,this,[],27),f=51;else if(f==53)E=J,I(this,373).length=S.shift(),I(this,76).length=S.shift(),k(68,this).length=S.shift(),k(40,this).length=S.shift(),I(this,254).length=S.shift(),m(this,268)[0]=S.shift(),k(314,this).length=S.shift(),k(230,this).length=S.shift(),Di=E,wZ=14,f=15;else if(f==30)T=62,h(),f=48;else if(f==74)x[HK++]=-~p+(~p^255)+(~p&255),p>>=8,f=68;else if(f==92)f=wZ!==undefined?15:77;else if(f==82)f=R==T$?2:67;else if(f==57)f=p>255?74:68;else{if(f==14)return Di;if(f==6)T=78,z=I(this,18),z.length>0&&y9(2,P(2,z.length).concat(z),373,this,15),C(373,this,P(1,this.K+1>>1),104),C(373,this,P(1,this[Sz].length)),n=this.xB?I(this,254):m(this,40),n.length>0&&y9(2,P(2,n.length).concat(n),230,this,127),O=I(this,230),O.length>4&&C(373,this,P(2,O.length).concat(O),126),X=0,X-=(k(373,this).length|0)+5,w=k(76,this),X+=(c=m(this,185),(c|2047)-~(c&2047)+-2048-(c&-2048)),w.length>4&&(X-=(w.length|0)+3),X>0&&C(373,this,P(2,X).concat(aZ(X)),10),f=22;else if(f==86)SF(490,D[1],244,D[2],this),f=15;else if(f==16)f=26;else if(f==59)f=w.length>1E6?45:51;else if(f==76)T=3,vK=atob(q),V=HK=0,x=[],f=87;else if(f==33)f=R==Sz?12:20;else if(f==97)D[1].push(m(this,373).length,I(this,76).length,k(68,this).length,k(40,this).length,I(this,254).length,k(268,this)[0],I(this,314).length,m(this,230).length),y(this,D[2],244),this.C[329]&&SF(490,m(this,329),244,8001,this),f=15;else if(f==98)f=V<vK.length?47:85;else if(f==17)b++,f=52;else if(f==91)f=R==ll?97:33;else if(f==19)U=a[b][this.oM](16),U.length==1&&(U="0"+U),J+=U,f=17;else if(f==46)q=D[1],f=76;else if(f==48)Z=K.next(),f=26;else if(f==2)Di=SF(490,D[1],244,8001,this),wZ=90,f=15;else if(f==88)J="!"+J,f=53;else if(f==49)T=40,this.T=R_,f=92;else if(f==47)p=vK.charCodeAt(V),f=57;else if(f==13)b=0,J="",f=56;else if(f==12)S=D[2],G$=P(2,(m(this,373).length|0)+2),R_=this.T,this.T=this,f=6;else if(f==8)H=Q,Q=u,f=7;else if(f==68)x[HK++]=p,f=73;else if(f==85)this.ra=x,this.G=this.ra.length<<3,B(274,[0,0,0],this),f=38;else if(f==15)T=41,Q=H,f=24;else if(f==56)f=52;else if(f==34)T=40,Gu(17,N,this,268),wZ=80,f=15;else if(f==83)Y.length=0,f=15;else if(f==99)T=40,f=48;else if(f==65){if(ME=(Y=m(this,302),typeof Symbol!="undefined"&&Symbol.iterator)&&Y[Symbol.iterator])d=ME.call(Y);else if(typeof Y.length=="number")d={next:l(0,Y,8)};else throw Error(String(Y)+" is not an iterable or ArrayLike");K=d,Z=K.next(),f=16}else if(f==73)V++,f=98;else if(f==43)throw cG;}}}catch(ba){if(cG=ba,T==41)throw ba;T==40?(wZ=43,f=15):T==62?(nD=ba,f=99):T==78?(wZ=43,f=49):T==3&&(N=ba,f=34)}}}}(),t.vm=0,t).sI=function(){return HG.call(this,24,8)},t).Sj=function(u,Q,D,Y,w){return QR.call(this,null,u,D,Y,17,Q,w)};var eF,Tu=(t.Nk=function(){return Cs.call(this,22,9)},g.prototype[kL]=[0,0,1,1,0,1,1],t.wp=0,/./),xF=ia.pop.bind(g.prototype[ll]),FM=function(u,Q){return(Q=On(11,16,75,9,"bg","error",null))&&u.eval(Q.createScript("1"))===1?function(D){return Q.createScript(D)}:function(D){return""+D}}(((eF=m6(40,(Tu[g.prototype.oM]=xF,g.prototype.A),{get:xF}),g).prototype.Z5=void 0,e));return(function(u){return g.prototype.Z5=u,p0});}).call(this);'].join('\n'))))(z)(Q.substr(0,v),Y,x,n,r,R,f),N[1]),g=N[0];break}else H==34?(K=22,h="FNL"+a,H=72):H==55&&(h="FNL"+z,H=50)}catch(m){if(K==22)throw m;K==75&&(a=m,H=34)}}}),V),[function(u){return g?g(u):"FNL~"},function(u){Z&&Z(u)}]};}).call(this);</script><div id="program" program-data="DfLEb//LsD6/ZaOHzev9RA4aWebX+QQKu/lPf6gmULhPd3O77pajI9MZ0+7jhumZZeE67Os4EEyoQ+TbFhvUdBUNCK9YZUi7GjNa90oAUezYsIaefCutrb6Ru53TKIWbjE1FNiQuRednMNgiIsHggoSBG5Ws/qn6DhdmQemxxk3Gqg/q4vaEAsHIgI673Nj1sCy2KRPYmbVOJdvMRjPf7odHpRwd4bC0FbnthW6oOrYiAjLoiWFRv4zM2AuOUR4qQZ4PQ1kyQWJE46Nm4KvqBoSrTwXaOFXdIxd4LYLyzd09ZL6HPHbx38N0c3bY+ZELdMSoSIRKtoWG5bMCqV2WAGnBgXOsS9YCbAR3VwIas0qOn0xSgcWsN9xf2lPwLrMxpj9C8Okm+CUp1nseSMLd/CoAkiYpQKnbqfI4y5ukpyOEWWGLJbb4a5/c2n3cJmLIUuDEGcpx3+UJxqAJphZTOMM85JZxflA8NhLPxG4ykBorWBvT2sFL2Ps5x+le83rarjEjbsjOh7MhKNr9NwXkEF0xl7yFNjFXOKsuNqSQFExzf2LjJz4NyN08j8vE5IBWkBXtoOKF5sFfaoPO+R5KzpUVcC6azWskTNZLEbFqwuePubpYAEiRrufbNfWJtl6zJHnoF4Lmua2g3Lz9tUHrq0PIHPymR9iqejKeiJEvsK8E0DsaBNhXuCdsAO9eGM65Z1i0b41G4mYjUBJSOf5wmABoHcmrkI7IRiVCSSxcy9jgHbcmRv8JFbwR9R6JdSooxn8RDlv4ICDS9IoUZ1IraAHZ3WNeYoXS68Hs0lF7NGSFuZnTGa116o/uJdla4D6wXrjr3cl72Ro2CIuC41CmZ+lfXjpxhosAPKOUvYQANSw50G+SCIxYQ/pPPLkthEyXPTE2t7Og+RspB3zcpnbpLHdk41NJE0THHFSC+d0fG3x83ds8AknDf8DtDQq8PY/6B+AleVDyBbk+10o/ykAqRZXl8MzcX/NV2ycrf/M3rFTTz1Ky4AxsWF2fmzhqxp/8g9/TiloqYbLYbhlx7bJ4wzPHcKVesF0QKDweUC7VLfB31ju85O+4JnSXk7IWIsGyEe8PuVJnan8OThx2h3eTeg/o4h8H0ftOZgc4/mOQv1Oz4NdsiMTLpV4Y2nDjSeUabUkitKoFAjfceYpB8lHKBz8SdVi0h8Q+u24WB0copilYZ7waOUX8q4MgfQY/R/iZZ+cAHG9PfBOJvE4C5SIShHfwzNGgcfRXYoVSkR5zi6tN4e6txdjC16JiugbwoUW5tTlSuTQomzFTUfGmMoqdVy+EdbainE1mNKrGUeH5W8bN+NZMGOyPQ3BmoBks4lRM+/dnfamFClwQSuwsaFMlqGeUqMPS/cyiBnTg6ddWpuvGfTQ3tSAbOIWdc4PrlUkHvpIn3gN0nP/nkB2DcRKS3LZ9I7yp5mQINyG4pXi3Nb13zmmuI6gY7hYQWWL/TfoGxdMu/4OnJRa5YmP7OivtLLAJvrwGygBixQ+ne6pwpss2goi2y9/fh2dJH+d7EgwRwTnmGOSuuuI10gNfPxIwda2KiCDDIc0oE/q5oizO+Xc4aqCrsWva5TGk5ou7V/tbrwM8uPKIF/6S8ge48zQ3pbGIsSc5iYueEqA3nOu3MOOPYAS5Qvv3fQAo1as/TJG9qnoykAjfmurUrRf4MSX1tc3ERPYvr0zo28B64NoF0j9NrkV69oJ8eJb7qRoJqszNPZjuvyAiN2T9XC6MDht4tHr4mkJcD+QohzEdCJg/lZZ58s74maR1eaCrCCEr2exK6Qns/HK2+gE+syqQOgYr1R+ec/D7sMQ1jk2/YQPa5pI3UU5nsb3ih7shtf9u6kZaFmT+8NyrdFBohQUGuHLlPxjD+GWaxMHcpngbnmYSKK4pjgEI18Pd3WQJw9jryXQGnPOg8Tuw+50Pq8lo2B+lRGAmEGfHaqAEPd0spgOccFwN3N0RoGghldt29QcBrY83IR/VOKv+Y0n2Qzm0SIJt7zY4NNbMLbO4rGg+0Vk8gk+L+ZEa1shvg2lo+fDj7V8wVjQfIYvyK/EoD7j+1AKI3UOSXdD7oS5suT9QlD9A+vQOx8XGJlx+kAc1UqJ/fIdLgu0mUTxKE8XneUGLv/+aldPonYYo0E2pQ90M0Wc/EFOvHL2bD3PUl8IURfND8rng12tdsI0+Uw4IyDQudIvoCz52G/0I4X8Jd3KpIYLXC07Dx7NCiHZti1yX229UX1R52yfyD2+GKFYRHlUTIZdlDZVP5SQZ8EyzUmyzAZO6Zd5WBkRhyOMyJKv9Jm3h+7pAQu9uNS5vkIox47KGDbBZncOZ/Vor235Q8zsF/2rdPerqVtkuY7IT0QOlOaHcX+4ZFopyoupaaiICXf8XwJVBjUyCh+9RtjPxMxkeVmRIs6f9igjTPCUbN5gHSILK6Wow0EgMRWwFWDiHfeuRcEyLLBm26+cDkVVO59g8361NzDSlgs83TTqLvnKj34zHta3/+MhUYXsLJzOd2qZ0WOc5Ne+jw1FO1ruCHF2tlrhA/NHuWE93wc6QMlYbq8ExPHlPuGSkl7IfJe3Tt3Tra8n4HXCJd/hBAzRqPHNEanxlgIn06h7UVa8AoW3+GELB7A8jP8J6GtQi+A1yrhV/+p29Ff/tGJJEnEJLexNnr59sQHCtBtCf3CmG2qiwDHqgFzUH4XFbsxnXkELsDuIssFGtbF/Pk3aJ0/UAaPuCJYN3XYsHr7MUtFho9vutpf1zWyIu8oSisMUQ0LmGcceFx98Zci/5V0avmug8X7Hez5/7XfGh1G9Yfk5bj2Byl22bkN/hluh8yxwFjgupnVFeCz+Z9PljFb/ieIsv13JvWvprZeF2dInfsg1OwYkdlwOZHql4+4xia7rSpNfAFyg+/UcjumDb+Uzphkiak/zvg/k/dOxOxZfpZJmbG3q05i1WG2E4i+1Ujqc88ebiSuCY/v0CRndr0qxOxJir2yI4GrqxRFo2ilGC60iwa3psLswsOk1NCMWPRVeOST1q6Nf95LCn/vAUpVmQ9X4e31q4M4KHP43oNrk+WcwpE8+d7U40c83zAIHzJGQHUuVj65sGXbWMhEszl+H8eFpM9q8FwWcxPayIYhhs+ImN1W2zwEe9TQxCfF5wEfO/Tc+tMJ9UCC4h8HkKVl8QPFBTPv6dHX7h95Pjgmndr+Fke3lQaUeHEVRiQXvHYfkUSWXd7ciZXnipOovVOg78zSHnlpXuprC+GmPfvdKNkTdlk/q2zvx+eteK6U8gP3tefcu9U/5OagN7yIEekbQXGeY7kEl1HvemoxMdz8PWow+wQ0yqLXPYGdf28FI62osRTLiIvemxFwd94137zGZQcwqR5whG3URBoTC8bjJtXF/mX2NXhZQGYV1Wj019pQtIeVNSG7bM+llzlWEnU8dZBz+fuNR8nQBoLwDX2a9IpM3tvUIq8R3S5obsV3rkqdtB2cG/hJoSySR0FVemEULDsqoRHGbYzgdREYDiuSFPtZ3kpP4zHSfEaqzxp/K4RlVCN4PgdmxPYbpbvHEWuj3IK6MTwqEiYCaNVq2Uj8cbVcUX1QLrXZq18mN1zrKv6tr8VqHM+iyJLSL47qvRqrjM3FvOgpSy813QtZf4mF+37Z2k4YcQgyXDdI6drqHpjvEIneAUy0sGgwe9KF9n/8Pe+PVNTrxt5nwHz9o75p7A+BirdiztvcwEnMYIfMogSJC0I0IG0hpLvtKEM2xA7q3jVTfIYoxHIak/7PL2j8zaKARmbDh9HBn76v0Vzmf+gRt0W1xboH+INTmwylShMvyJXtwrubwVItsAeqg6Y82SgZwkzaGps6Gla52V8GCucy+iAi3XAXCtuUR9P3OCO9r3FedmQlDgYrzgPhg4QZsReVMYrF8Mx/GyPhbQ/KUPBcWAQsvcGXs0wRz+A2ZvQkEo1eiL8FUbDGViTelOCA36mhpmKefm2YZF6ocxmfF1DVdjEVttDdt8fLwpsTIdccPU1W1friEcS+1FSEwESHZfx3ZxARGikWfXA4x97r3Jiv2STswsVFeQ2Xh+BZbF/m8XsLRrQVdZHtGwsON8/O0Gji/1QSyc7wi56kVHCyRD6OA/Lv5z+krRDONSLMp/e9ziVEZxo6ZmpykQgF2DglH3YAJE1XV7wd7o9ou/vLkw4JSexr7KVP7oFPgg3oW4P1U6ovx3/93HCRdU8wIIdV5PKU97GRPHLJRHFr0NmEiL1FLGPR9vtA5jJBAj/WX02cLKzAnsAg+K4mdXOMxiUKIh0Ql3RMPzo1ziprChMyfJXhdT9TbL21OH9Limk4ABxHvfPd02ptgXXCgQJpX0mxyHlqY/7UmGc2rQ8/1ZfnhQ3OFh660vvO2bRVOEFszZ+d3EPvqXTI6zB0ZgfnIdAC+HW/sZcvI6dx78UvTldXUQiAdP5IEUCWOe27oI3IorlDmAreaCd0ZVtcT0WC272X7hct3HBhE5igMWFERttA6UFin7pKgpY4wNJd7pqXvuGWeaOeUbuitu7eVTzsBRmVn2hMKCHsN7nDt87XjiH2O6LP0UM8Zb8zXajVWB8ZQUD0XJji/1IypL752UabD1CAwfKVtGUXrJrzjry6HxolSEuboZLyFkJSgNfHny5Ps1E9qG3U6uL/bBtp2nDV8eGRY2/KtjSUmXM7ZgikDYDAbre+xe6rE7wYPlT1h2tqD5tumz2kMEitoGByKzPF1Ph2ZWcraYRLdUStIyD/l/B1Jph+w/9u2XVQBMjSmF5YyWhKaEb7v/9xIbXUPnrapUkWlgwZzZlITFRJoIcPwXx5nVtudohDmJhXejCw+IeYhKF0Da9RJjedmM413OKCXhRypqUaERroqakD4atLyC0yBq+ciem8CLTcLxI32zpEgMxf+Pr05D7/ziEiOJ8ghD9LITVnsuWLv/M0AbozmyS1jk/v19FXcPDmhB6xm4vITBkiF88eBc1QlqBxCpLvy0FNt9zYIrTSuptNhW8p3Xcnzqlfm7rlZfFpxf8vNHlggihVHIS/vJ05Jy8jv1m9CYnOme4UAV96MXOVvaAwaoLqN0bOyPLJB2+z5gs0dOElozWfPwhydAioJBeCHGs4qms6cSolslfnP/REwaNccrZA8oS8/t+LcaySOh5Xnx/08ogzigd+uck0a8uN1xVWKanSQlN0VJztZZYbCCPoeUrMiAJQodAcYaL0IvpIIzLNWTD5NCBiG8PHLCEGgM6Y9XjWK/qhds5ffzEzt7j1LUwrh3UKzqOeR+Lzhp7JpnjFBxS0ESY9MrXfMtvBLjVHvI29d1ZbwsFOWkiXoMNK3MgzLQfEdJBjev+KPjgpykion9av5lceHzWqlR1bDKMxJuWUNUCgZvtE9RXRcI8r+XBv3GlmhE3ZfWQlGubS1eOsI95igoWYeR9N3RCM3J8ZXZPZ1jnV0OkSLpgRm9S/UjvbbdSnoG1ez+chAN/9P21tNgdV0O8G2KamFyI5t03LmMTJo0zMCoVFaF92hqcrbEhbHJXbW4QS+0CVSBuqtVU+wU1FFd22wRW9chA35NxV7ix3HO6YIceFSFfBi+FRQwQDIt/85NZDR8NojEvabF4/QloIcZjcGyB8tMHmiPiz20FgXvtMoAU1NeL2G8weqoGWbcUYYy3qx7ypeWyXhlVcbA1YaOmfqEgZlif2L7ZQQDOxdmTXC5hF/T0ObLCCLR4IpNQO6wL/LlVQwIpOoeuNWXXKyIClp53ZUnAP9fqrIfPfbLKowo/fLSo49P4WWMFwPBIXsTSQPineQTOm5jOK22bWPPqBuMOBYW+BQKdU0Nytd92Yxy0LucV9fsjb48f+8KQw59XaCVaXMMs4DWmuTendhU0v2SzSQycbWoJh2jQMAT2Bqv4RjzrjxoaOKRUUhpUnUDlZQBkTHDsDhLzz7vjuOGlqxe5TA5Gm5+nulY6VdQaotkuObJ1uIwD6naLSwPMbYz3WG2BFPcDwEnLgczFxx2cQKdObFEpyxvjwLbngh+hORbbnhFV9TK2unzyZKZOO9/PySCI8hnZHgciO3XAC6ae8Kvx8vBScVACkt094AvlOQ+mUCXXOn0Af9MAFdDkVB/CAesMfNtgM5C99Jl6X3x14Yea4R3b6Zn12cICdsBLX34vUrQdA5dyWRS+inb0LFnFsgbMnq9RdGCWmOcolE0aIhkpPp+aYub9ilCjUUgsGObN/vngTppcOolo2Kxfi2qt2KKtnl+F1hstCJpsNYd1UQfIA8AEQ3ewuRDzLb+0zYAYiGudV8ALx5V+EEH4ywHRyV4WADF9IJu9SLjxGNp7HYoNMioznLSF2Ms8RNT2baS6ZyRtJidCuF4zE/HJlgd0WYUKgdsUcPeMLOYvnfTYOFF9keMve3C6EkX/PoWmJ/mqld+qWc9+2Bml6Pg56iH48rv9eJREnI1Ys5XxbXfQx+U38Ez9eMJgz+01eiFasC58a2Z5s3ky+2nv9fr+Qq5sj3DAl1LuietQhGyjtOCfqx68HLq8QZH0WZyjxgOGQqnx3l96Aor8JGkOT+Pvv5vZnXgsHiHty8mGadVIDPT9SAMUqHVeKPK+IG3sRNsIcfokar8lEF7rKHXPeB4CYxQS+JvhZbxDuo+K4tX0FqBlnDW74qh4mHleK6JyEvUSmc3bW5jtT1a7nL6n9PtbNwBlqYSdrLKq3CDHgkAQ7VRMiAlzd4pXDDiJ9YPN2nZNV8De5byQkstcFCaDqrdvMPlYg6d+8GmP61C/cjNtXMm8SoI83C81nUtULNwXWW0E4dVrPLeLv6WoMgulAJmktWdTutt5EinlXzQgYYYRr1L0W1a7qMDFOdrW2CiICgEIzIlK3VkMjf6xcWNhfo+5IOHp5bQ8+MI62r8Qm6wdB06hzf5gLSR1/kMJcSoH+XC6DMf0UPip77YmsgKOGlV9lNA5rqdKsSzy38zG8reYhaY8NhUPDeRt2ofyjMX/4WKOPbiWAVIY1BTl9rvgpyz+mPWVXxc2TQn0v2WJYg/VYQNGI9JXE0WneY0YKnwR/GI5IqhKuDqkMuPT6cHblgHJLIjcrcS7rdKGUFbujkDoX3izqrvpJ/vFg93b/drK717Puo7UWjzY3xS/2ZXQ371aL0EoT4uleo7ZMf0LGsgmbW8smW8kBZevUtAJv6NZeNzHH5+bFkHsjSKGUgnCCVCJyyCF2d3h1fWt6Aq60/HliCbf8bGisiC3qsdpeGbiOyWzfpFFnfilbyOpLCFqm4Pf+JlDLCgGwupJR0IuRjfCI7XMlEb3RuuvmjKNYYCvI75KeZYAnTsBzKWToLcp6AZxLhdZHE6uBrhFlZ8Q9N5J5QwRW9Zq9nnXLZ2HJ6wYtXF81Gi2PK/kCAOzbj2ECw/WP7hFmajydTtwAa+SnvEemLsdys/c+R8AKCiuFB1JJI8lyvy4Q+ibju1TQlRfVDmBurp5Z0p6ErRDRSRyxB0q/g1BAIJDngnn/i42jhcffy0Qu9SYBo7WksSD+q+sdbmI7SyYQu/n7FgdqMGuYk3aFOHWsVdBdDadu4R+8QjL0llJXgLu9DIysJ/H3uRJGXanUbNKUTM7R6rLXqUeHBUeSz75Ful6bH+FpdMRD1z7yc/1HMmfW6xUCPM85Y/0GNZemkrZWeYjO23L3ppWsdDlXgs5QqZmXUnPItNui13mdgH9SW7U8i3DwQMXhX5qe3ltdCDE3UsTahGwfumxJtqhaXeI2jCHY58rbA823aeVm5/VH6O6eCS37au6GREaiVjx2r911kr8TSVjvcCflb2Gpv2BMc2vCskXUU/Nw7XmVqZDuYziqIuO4CmCvBp/EUtOaB/rRxP/kbVxSlq7hO4L9bSi+/6MvPB08ZxlyiQMo8lZQigwK4K9EdSY+bphTfygtkhg8l28wuGZT2bsHzV+FIqfycPBGWj9bkxtQcutbfk8MUXSqFBuMjtbWd2dZR36ibx738t/2kFeMWEXp50FS5T9x0I3kr8s4jeGurFye2ra/6qc8TqhaPUB2O9UytcAATVFIxDe6rKfrahdngh1P407enFehkaGpgTu+GlTUV7Tw+86o99hX10uj0mPqvTMCgq1zIawNnlIfx8Oul6fP4lPhStXfn/1OQsA/mZttD0B6khnubMFgEgWiQy3RQqi6OblEhmvAd7o1eLqDWI36j8Ogo4HsZARbbnoHPVewq9cl3xULorPaElTKyQxgWEA3+5ynn+r3aZbdykGxlyg5jo1zweTlrF2VUeoCku8KvBkjDZLIK8C5/uyaZHF6CoqBQ6vd6lC5W6w0R8lEWsOCDFwT4/SFdtCf0nYZ1TaJSOQwkDxbaT27Cf+MKZ4R40YZz51ANwkzBaaVXMc+ptG2/ZzK8ifFe548LNpjffJwb+Q9kbPl/WHfv+9VtS1wvRuycXjOiSAnxL6o6ulmWVA1NWJxRLjgJcgydNP5BldIYCchny4h3USYKAmCAKRtSkKCoE7lBXuFO4ETBAK27Ip/ZqEOi6X0FgdHIFyXSkmM8BGcylF7OLxTyKloZKFrw35xKU/JP/dN4YNRF3XbH1LESZoyCSOFqqqcwGOOGRvm6h9CEy1VT2ji2YfBXSW2GVWOLxDnZK6TzBrPphqKuW42HHo7binlw9Qa+aFtz9oEn7SmmNeLoI5hYQIPkFOsSatym6397/FMeqI3QcB0OIwKT+CxC2vHAEDh2F9dzLeFoYQNvl/xOrf0xoeJ8D6BIcySufEClDirFQnNY3sDGSsiUyqhugXFXCJA75BGAG9yCUScIlHd5a7xi0Pwf7ep1pXjowkP3wyqa9PXANMKAo4OJV+9d7QpOqB3J88RT/uluZiPxkpdRh4i3yrs7NZ+espp8vcee8HYyDclne+aHPMbfjky5SEuIS05SnjXzdGCeouIGryZQg1VyqBv0pJfsc0s4yZFEJGtgoFTEmpm4HYSq7ixYOaq05bByEJCdOTRc5GMk+ZF0V/Xb/UrKMGC5mD9jiZnGdElL6DEZnlQoY+EVYPqcxpovEFWVfMxeBV7SJL/n8/SmzQ0EHoyG9P6GLjSO6Gs4pSA+U7L/4OaNkXOq3dsstU0rHoVUtclDfKqYVg03GWHJsObew5DxmAHcvNdz+VCbnuQzv7rjtZzEPgzjPvx/rFesBmJLQ8+npdmlGFU+Ceo/LysOEiMQ5pCKvBtj6xBBDStMhcsS4Phh7jshvFJGuJbr+/0vFi35UZGvRIiDzU7d9cl0xuXDMzKKNTDx8gJyy4MbL3CyPgwVqwdsk64MRNBDsmJqP6HQPNckZTZRmS7SqbdysXl/Qpr+6/owuo4xZYFGFavnoWeMVQzGjT1E3OVpMCP7NEWh5jAwQU75bKYH4NFaKHtCrkVuZsnPSpXzO7JAie06s2D1cL6QS4wInsX60q+pjjfUCNsUzdh93maSq+vUyoNhketxgnEkNGn+xkmYLHSqV6QUJPHVe3j+2YWm1YLGcqF45N9nNB81xy6faeVjWIm1y3JRFzMQ4bZw3Qot5J6a92JONc4sacYFTf8fxET6LW+TNGagRuUSVpQTZ23aX+2Jmw21SXAVoXPuOG2JdWW9AIHnnNbwQ5eOdW8Oeml74HHkibsTXyajdbJBZT5RUydEih/4FZZRkP+HtgYEL5qJVBrWJiH8YVHlvAMpVwpWA2A1tXcBZBRyJauGepk1qlfP0CMXoLwrr4zrrCGcZiTY7/hJAmbyyr/OS2UAiEIPpMwSbnFrsR1u9cGJgbUDwPCDsIWdEDYFwmMuTvbGrqSzJfAGc2+Mcpf+Qr7zPSge2B9Jgb8y6CZxN3w71QBnBCHUnwojqvIA5/PJ2JzJh12YrhAqG0duU2edXKCJfllTROkhZ1xwWGY76T55sCxM4uzJCBM/gJFUWBKC76qbDPVEmtNFjQl6T2J4v1RmnrhXxadv1m4ubDAMZnmqQvMbEIMC35uaiybLwOAGgNVAxw0T2N5vww6Qd8p/ozjwnPHl5xmeaI2DmJ2j6GqVXBomnoA6wPZTyrLCgTNoNgn1hafDqag31XBk6PT8xx/UOPeN97wjH0utD5twsgxdVMiOuLyQSEEi12zkfNQIAV07pHbobXnI55/WDgghPjUu/VQWQuwkcIFSijgbOVSiRQoIPk6ZW3m7i2Ilu8gNyrOyFB6VZ0aNgCiybO7AqScit+agVSGPbzuY/MuTtax93YAH+WdYxzMnqvT1YR5bfrFmiOFyJGlBiNcDi0KrCn/NFcVBGR7obpykPN2bFRTLnms5yUjAdZ1XEjpCgUT6MKgfBhtFsYFrnIkWlsrnS/tDS6kGnEydU9LowRqBIAZ9B7V4wvYpYqqXG6sQHc+sp7HJfmZqQjCfsGC4OxObr1PztvCv8bItHRCrk+CDxZ+39rtvQYAh3+mb2KIAvrzdH4F7vL1o5bwW+wlF19OUfUvFG/g2HF3Veb8BThxeJy/K9PUN/8EDrizaAmahBod7TdOFOteYzvBSqcllrEhvouMQ8kD5oYFLfMSWWKS7xcuYXAohI+HiMoShzohHA9I7qmV5szVL8re2p2HEpMU3LeJWXty0jI4R4fSoA7YMkfYlbiVdkthN1T3ZBulllQM/700kyn2rE4kXe3L/WFH9uLe2uUj/lFdpKKXi4mkus4h9dPGb24QxdAgveAMAjZ4aTVWz6AXuw/cjTtXSscK+FDjI4kkV5WMes85S0b/hgK59XSGFqAIRcAVrN47UxjamW4OVtFvClR1CAlPoNIVVwuQ2FovFbLLyh33A3UeIo4a9k+M0V1EUkCh6MEc+VxtE7+/cX6FlrYnc9TfK9m4FoBEbDzNR8IQZlC6C/nrMOt2qChVYeAAO67mhd5Yjx9impdB8VQH59yc/7I2e+ozY6SGLQbRJUukLd6MaAzKYdEc6XnAVCZr3koA0dcG3PaczOOFcAjkUDezPttoffQeJUn0yVH7TbPIgc2XZzLXBKfXE3RdripAS+Gf3/7CaZU4xiEbKswrSega68FoiPI70WdzK4jwbCAaCbWxE7pCvvepjSBIRhHxYfdIrWa8Yul5O+kj8K5CAGJ/W+eV8yDQXTGMH6J46aLAAoEp9uv3VGi8a2ud7f+iiM18971BjC6hFXZWxVm/skFVrF0nzBNBa80eU+mN53YwYGBqj0fNjSnn+evuwePWyQp4Ye7Zmzzwwzx2HVsla9gDzouUqN8iRzLhfNjoatJQOYAYP0BYcW2zKDBr2Zb7cs/trfNAb6KWkh7oASh+iIsmaSyfBKPxoddEw3J2HsVTCz8AGmq5UbFXm+P9F3D3yDm/NQWN19LapU8Ry0iCwjbErewahlOcG5GsIDC6XPHuOo6+egFP3bGNLJat53Blt1nVHV4uXEbJT4EGbPIkSkfEcqOqRebQDd/1shZPVJo7O4I4WRdCB81tWn5pHqmeKRs6yHcot6B4fsD61JiIqjBWkXY7BnB+k6cvQkryKolX6oYRNse9JfVJ01qVOWX7jHwepd9IWziU0vdPyzHK5pXQq9E/LOm4gF3LvxNReH7h/kQQp36VkLisL9Lb8ZNglkQHwx+kJTxQgPlN8ZMwqs/c43A0K05ETstQqgAm7yGA1ZuCe95D/WhIZLDdnLe6kWmWG2oZY5CSdA32CNvakXe3Q2BycpKCkVbFAQTR0IPjwgrItfuJU0A8wiktGrGoiVomjplGjZev43GsZ2izlwOCV9LQjmbDsDTl1pz7fozqYAUaTvQwCri1kTvKfNlayJOCJ6jk1qckCDWQsewitEisBteFHsaOF6yRWeNwYKoYFccStg7fCJb/mixDAUheqetuZy1v4Ocmjd2AaDxjd4jYIGkoWVWhiSXZm+O6c26wUihoSpvczv4kF95zBcJs6bfRxYCnPRWGLEJhM2T6Jl16b4ulvPyzut0gmjuPsQ09DLF/iLFShiOnv+9sm1fTG62rnkwqYYPs4AR9BbzlI9qEcV4Ko/ZkhwgP32dxF0x9Row7EOIJYPKPHzuyrKCR3Xh/Kf7/OuvB3BhvZ0cl1i6sWXxCIFsShyWZUb3GUO+u0cexmYNbDnHz5oDy1aJRxUGeEmwDE1GjMSOgcQb8almGHSWOaXUj1Gu76PbMXD6D2pJORLlDvCgCemGGx648SJwLyqyH2YqjoLQR9o9hunTw+FWfu96kVN700Uh8eJOIXujvCzUK7Be1I9UhEWhTn1u1NN6COac/UC65OqFNBOd7PXIkKANgSbBDo4KaOSvC02+d/lxaZH56pAY7jdi+MuhtX/u2Gud7dGnRMc5ZjaCSmjHc44MjIKwhCm8jJ60m4m866ZNkfIAOKKD7iaEoWaL9xGytlJTwR1pRk1jICUkqyFHgXEjtzRIcnoTS6/Dzt8SfCungUNqYWxrgHe6BjQaM/NMb6Ndx+Tza5hDvXQGp2bJv+A+/9B+2FAT1IWJ+xSVwL59UGdUty2JBRB6cIFbVjxkDNMgCgJpIepbn7soelUXZZk9upBIMZ6cadiAL/4Zj9mqMyTRD2uZ4c5Yk5EVyzMZkFzxkSfo1tBUVRgc4c/JciZtWyBp8kjBp0R01eBqUEdsGww8JOJyYhM3GyhsF0ww4fyDXZ/4K1ko5vyZh/D1SKk/fW+l1HCZ8H/h0a50aazpBPiKekPXaX1KtWiHtLp4MROASqnx/IydueXWdJ4iBmVXhCK3W2dBXeJ3DRh8ykogiIUdg0OBDR2vwTBcnBn3Up7jA7jiaSr7vJ5r99utBSyH1gx6qzCgIrPKsmKvGxAPac22YYO0KeRxDEYz/uJqO1uBcLdc0OuFTazfRwot6VJWuQbd7+nIsFnI/YRM0E5ccQXgYjyanC1mYb30SCKW1X8pWvnLdwCjRsGEvgb3kdMy8Ler96hbBD2fQd3U6MCEAh+Ds5r2kRmHuU3ZgSHI58QJYjVk5LZjkFD4D+xx29Wjl5OsE++FbnoPPHD2Uil+R1mKCFo6OvblfrY7ny8kc4PDsMf7mUrd+wuKEH20zlQvYZsEpBFB/mNtIve3k1rbMAvcQql6Cj5Oow01nLZYzM0drru4AlSgCIJek3AP4SbW1QzN0rUB+p43t3jcizbIAErdkIEyckKwPGebJDaiUkzlOQrYznAHwMxR2UsLJidM8cfZ9TNsO/ySSHj8IbLWEgX6KFNQyH5FP1A7ygBFapKakOp3id7tcXNFx3B2eK+u5N8ppW9+F5KyJ1C5YMMeueu2bN7jQfxY+w7YxFWg+9j0qKUJ3GMMAhyOs9eMWdLKFYfnug63tJEtJjhFCqV1qv1bdwNFVa+cmkd518ANv+YLd6kU61fgiM67ittaNtFlVDE29QGYEAAv1yKn0GIu/VGQx97DnR4y44ZrMzyFsLqAMEdqKPn0g8+Z/M9UcPHgzWCS8sg0hoGDmDGi4s/M+ni3H/9JYrO2u/bQN11d9+xAfrCNo6wCxZPsBlokFkUzTYcporrbYbE/f/uJPCDqtlb9GrhK3/naHxWFN/Xau7GRln/0xnHnmKkuVxpQeWt/MF0GzpqkyojaseSGMEEbps1twNJMwssMHbAkfGrl2s89Xd9oUG/S5CRy5WrSdKLpa2eYu7WnX62ueYeFJzO7liVCFbLrEsu4G0hC3k1LwZb8CW31zkgi/8r+IDnhGRAx6Wibx6QDHDah+C3kjC7LsUt4vAU46XnxunGpaF1gtXPE8RO/g3vGJnT8VK5q0vkPaYZ7/EFQQ9UrGBiX/C4b17yZCjJR2bn8NIyrwBgbvJJ30JBevYOi/AUnNOeshI3qqfiD7EXXKiqAsYNs3HWPLljm9Hz0y6w/XWPNzoTAfhXE9iZjXpU3Zmrfw9J+41BxBW9VhvWTfDV99IJPh0rAqSVpbNfnCieTKYmM9nwh6unLVh8F8YZKv5Cze0mfvKAIg8Zv7B+Y3KITzDY3kAgHuzgUnJ6BTY4KUouMe/asQoqaFdADIz5zX0+tilWiqq5d0IuT6CN0j6qSVsielnrAj298nTn3VLUgh4Ndu6BSLL1/5zfFOrBGw+9tTW7y4OnWMdxml9PozEjDcGOJ2yLHvwVobxFCUr6LUZXlglmMhlTTqnaNh0tbDagCe5P+Cfx6fjLMtn+sFTZ2ryFVZG2uvoQ9w7HZegWoVkG6vaBDgfHz7vFxDBjSIbQJrepzX86hu3TTeJmA6hqde11dByygf+VukbMHWzOTjVSew4V0Z/z7cFBOhUmaRA9hQtg4ZAk2ppZYZdf3sO4+Jbfe7SiTSlUdDweQzPAwB+PRRLywvKy09Dy5buan0nJ8DalJBRJPeftp/J8SHUZeNe4lCriXdSdLpTcpMdnvGkoJjSSq3rXDYb/4Vo11HsTi4KHgAXuoqmP1y9XgpWz4Cnc+ZFEkhzeQ6OSSIJvdz/yHS9iOBaOxg7JlfWEhkAppdJrWIoQ5CdLBGNZW8wxy63gL5Wn3kGZt0IaYVYQPWybCodLIXz3P6d9021Dsj8YrzjHLZ+HkCApNeFlwRHrw4bBQngtxZQe4ahkyq0e2CeN/qr0OyAwdzLHd+yjpZc3Cp6EGuh8Bey1oiUtZOaPDJMZwPS7ucPtZYlvyVbJQsBS7uVT7OHyGCFsN36n71NLAhlUd4zHLQrO7XQQdAyQ8EzIwgGz7j6XAPUnsO7JHvxpmPPxuEkgr1UxfBPj0SE7Vysluf4PgZkK5tQbVjOz65wdt+2EWAHWFoYBoGRX0TzOo8OSu6+1AVPMdrJms/8y+X/VmUwjPjpkK87XvNobctL8VydnEROZckl4ReM8sRACDNJtQtK1umOj1kQ9k06rCOKjUT7dFXik62w9wvDNzhKo+So/un0wn2+EkpRMgnt3yXH/5Ps22oV9iLfUFr0BIMLeUMp/ETQg2prXh10mj0GP1r0TdUJjNlgci7qR6RdXi835CtS5+nfhrA5f1cUO8Gt+dG7BcExdu6sly+Nupr+r5vdAP/eovhg7wjDDO+W2cOGgtMQ7TK2nW0uEDY1SLqOo/Bhr291M5yRZuZI3pls8vPK+DIMrvVweF7ySwLL437TF4HQrb9NqSuoDVjH3S8Z675A3626WXPCn8qpF5BKHbxK2ESUV4Gi/7cSwEtf98ssZjLACvxRQn3StrUqn1WWLi9Hs75XbgroJTB5Qb0HRRtTY/oyyIG7lOrVzlhr0pszjvV1wFUPQx5BAAuMyvOJQptqxfGHvRI3kNap0r+fGfjIOnGPFO6w1+rWlWZwjXwGoUY1HeiUo9rHUc2Y6xGN/ilK/0wt0gBs8IW8fcSWTlo83c8ijmrbSQPWRp4ppWxmiC7PDiyocNQcVoqiD7J3X/ztfxc1McNdj7TzEjMuOJVHI9440FQLL/d532arnmvIdpbvOmJK5Z4V6k5ILzi19Ngl50Ajwp6o0jGnLy2hFUSkciR/HosHhsyNceHA+Q5HxIhaQVw2afBL/UHQQIhq7/MtW6tMZIT1i1JZ6X1C1SE5OMrhN3LpqMnVW8kk9Ft6gdAMu60W7WjVAIYUDNDuXqIOvPCyVqblCoK+oWPPk3bD3G2tlmoznIP3U2Qo88Yap7a3NdUC1M8M/YMKA917NNpwDWT0oJiS7bIKX4F6soTN97Jn4/PL/kfjsVMS0hdBrBneUzQqgC1A3sndNz5f4tafKi4LUEAqVGeMT8xL8yDb6X0Wa+YLeFSXyLgKI6ski1zqF1ZN5628xBa6hziHH6eIoBQSN98K4ucXeEXDE2hFp9GviXX8m5Nio9MmI0FfjyMG/7a8p6t9XnBXHscMeYd3yLmhkrfX/U02wkCuo3dCQlckUDUAB4DaKqgDnEQlVkl667u03cLPhN2+sUMeQRVObft6kYOVlFE6mMUXKQedfxz6r6XSGuC95fypdMK0q4nDR6gQD6huJTU4pGBEFcXitrH/6c0NeRUsJn5fj0YnJJjJOd0DWyEoAjKs3pHkJ+H3ulHGsUMGsth24xLuTPnxZzJ3eosJOgYyqcIzgrM8kfsnpWnJ5T8RLqgF5o0kGSsxoE6M5yS4ZdIOKvsxcRsrzVmyJdKSQcNZqNB2nB6SknyFShnKbkDIgLlML886fJexhtvtKt5+zyXhBwgtVK6RtGmHEPtA+hkX3N+kMzldpAwiU4BD2o+RQjkz6Zm/mYFJ3I9L8WgLKwPqryuh8kLFhjZ1T4CbLUZzR1B4pduUB54ewV6bdvY9BsB3jmqLyn3PFjGHZybV1n1JSwaZhCdCfZqBcCpsPfVtWDCIN3g2YpdiTkD448BCJV8+I5Xp+GO+TfGE/IlRpNUegiiRSN8KAODClyizNBGkhPe+bVPiZKyV7pXNRxn3IjTiw2QKJaY98mf7ShZ8zS5XZobgZC7DsC89yqFG3LrxxKuoCtTHCDHEjEFvGygZtM/Sep7xfW5OifpAlRtMABJhdHe0+JdAVa6qBq/1jEGmcI06JYIRI6qrCKFdPswI9bz5CzhLAX+fltdv6CxvPq8/Vh9rsUntDha6GzeZUEaUUAAY0orjko3kpzo/zWDlBAIbv12tj6RrlOttwZXNU/uQ/Kx2pGm+9bmHUxF2J/SeDh86xyLyyKBOGdqe0resO/KCeBd5kOSc6P94IkBuZp1Tdcwio/DKQ5GKAAA/9tT1dMauks+pCysev9g6FNAmfixPKVU3tzCqnfq+8M2kIJIFHII5g9q3gzB833WPXJGkLhrZVviuIc1d27Qg7uSZ9A2o0jnaEWl9/5Oub103Imp2R0/BRZRPMQga374vo4YoXLcM5elgiKmSEtObfqOTn+IlQW67Mi6GvDOJ1A1iZd+Gh7ug56QwLV0gR5fHX5ee6CmOd1jSHtftyWmvvilpCgXtPkr1Vqy8dnezRgOgWfjVS3fRoYiNyS8J613D+luyr+a/sQo5ag33IVpCYjQQal37i0FTD+oCcbcuT2i8nd3DiNDxVO7S78g7pjuq7YHLJvtySv+cPvPH7kJe7X5j4+KAyVi3DN9cOP8UqZPVzzj5kz9I6QiJW0lrxDt7jd2VXXosvZR6cJW2znp1mYb8gH3Xhi2nObriQHI5j1K6Rtg3JzoPL8pGDf4QOyySqb6Tgt5dQqjR4ridJlskKiKsfZjSXJhcFqohMDNCWH4kJiuh2UvEerfo8VFEBecTlmo57ySjWTimbqnm2P2IsugK5Y+0g/eDxCd5yo0M9hFU19pX/FxRO/CPt4bAsG05I+AKSkdOw+QL3TbkhMpaXupE3WyDoZvCoVTPIHrXPjrBj3t0yhyYIWr6B8Y4ZTOcDBuL0Lkvt2FVvDFk/OBTI9/TfIzMn5kZjdbu7kSDppNk8TCxgZQwRolui1VV5gaoDwR9tE0fZqK++Vr8zsdQ7c7UrJbY+MtB3qp+iZrVSI9r0k9ZP94y3qr2eWywJQLd5MvlAqSEGKAOa6oH+NB4iKFZzx3Sb6jqFWk3n6LNXUsZgw/+BgTayRPIunMxloIfJTAe/4CI+TQo6g7uCWgAYKyCuWSreAzyOeJHz6HjFi8vLavsZcn304/pr8TBcpD2Gysko22JpR3YZ3LGPfG/ulHivmfUz4JgLZK+egRMAMICygngMLBeGnUJjfW6N2Vc1lHW9ICi39ShMoFu/WiCzIE6LxHvS0UT/dVQTaecly1eRyKsflPmi9QvAoQHPBVeCvJn/w9zjhV0J9qWNpPtbliGmkhzzCK/t8cNCu9XjI3BY4svKZdoemMFy7ybOeJjTzd/PJzmsqE8Y0undvjvOYfyuLTlxukjXs11ZVGDSw1RLwXj/vJ1xiDoBxFqPNVkwR2bicc0tumVh7FSwK8v3pJEnB6gyutFgc5qbO31hUHE9EqJH7xCAMsjPVpbvh/VttEgnm5Vxg6p4233r55KhTsEeHGZElPnFDpYedOZHH+soISoheD7JRLrhzxsriBYZRLOT/TDiv4jQ/LYZUbRBwmNQvdmLrI7kKw1+CsM9n8DBBOpgj+LybkdiDK9Op56/5hwj0JLjDOEMYc1XQ8+dY1sX7/D1c2ZBSOfZ8L+HvsArdspzb6oD34mxnHYSS2DUTTwV2pjYzllqkcMMInueINOluZLKOmhRmSK8Rn4+tJgyTRLMWOEbAmmvVq7FlShkOMbcqK/1W99Cl5UeYikptvluLXwUOyOgNMYocoGcS1fWOqcDPnyt/l9NrMkZvaw6CT8QRv0hJmJdf/Kxo+OmDTr6c+L8HxUf2mmfTXQqdD1t4jrRZ9y8vSy6SMJAd+VoHK+2gU6YKQN0J452+CRYPEpIK9b6oSahlGyLEFCqhLTM2KAbg7VJ3i0zBYG1cDXEdrLEcRp1u5oScc3Zvy/nIzQzfO6lP92Ftk1Hbi5OJUxnrIWjhF+ILpKWJSr28EC3CbccY1+QABaN0tsYkxwKRfXKBZ1gaeiaxzqm8AsopQyQX4mfpJ0pirfjGTJi+OVwXydMB01ARhbwhZ/Y7Wtk5tXQbOUVx4m08kp8j1MvHHSN/9NkA52oLouXZ4B5OyyAUBVAdKfikukCOzw+ys+K5TzfoOOVItqBJC/6C5S5JnhG0Pa8RAQpMZH6SLWsWB2LE/SEKpMgr4WxsYEsuE2K1jkDn0+4O6yeVY19EkeqvtOCg3718zk68kdc64+mbkNiPrvLrgEq2eDGpECaoU65YhFLe2cutVNH7EQRfsYQGq8PLr2ldVGkZpAFoNzjrQ1iXIKqWVLCK2kuP7dE/+AwErfM/VOVRvemUR2l1sVLZdi3NAJwA2DIHUIuJu+uutROIhQDjOvfNl9YT2n8ZH3PreVxH4+9Bxi96myzDEMJHh6V6AhNmXyqVQX1V3yiMJ8NXAoN9r0ooRRA5cTXHC5y+aMmUBWgnVk/bD4NalEKqLhkAMHf7CcavmN0+zcXOoT7w9YOQTCGDzn3nnhsvHseATRddy5iJWeU8EHV/9E/HGBd6HpK4mWClG4HfcaUUwantHDTwEzqddXT+l9mqjySgTIcvSuvLW8ka6nNlmyi0q+MjLUqjJrxWFT3LKsf1mu4SmazzKlBrH/piTKcgp+WxA7FBFxpF5P3sseQLQkeSZs3OZ/D/PWPDGyuKVVLnLG0+Dcwo8rcOhbQfVqXwo3suhDCIvnmI7MB+/78GPiALxMCXX6/WcI6etXBdVkGROyQ2gO5iKPLsov6oOjMMRTF+9UtdR0FTDj0LgK8/TOjjEV4WXDJ/hcAH9zBHv3Rk1lQsMBt2qdMx9VxnIjuk0/SAqKzrL3Gyi+BS5C2EX+z+/AX8EebfqKzgGoBSzyF2M0wp+c2rfwtcLL1W/MuPaHeOL/qxvnX8oHYSc2Up8WBdIwnFbswTUSdyeEtHSfpICNdmSLiuIzqVEOHA9/AAe4LNHUCZpW7r480FDJiuzjmKMk286+LBUzck5i48BI5N/KvhqxAPdS0vOD41qklKxZ9uQIH9Z1/zA31ffUu12emBmieyW2+Fjt/liGNlIZiN4goy+hqs8pQTkbU1Bc4WJsj/fLaPqaiBuI7m4GiHVLeoSJx29jOq7gIrGPZ37YjQYFYQ1EaFzG06iXJH+BkC8T+3mbhZjIBeMRJLblpBalSmUOsZFufLki8tEmcqKCD8Y1bNrc2PP5H255w3CIBM5Q0hybiAjVhtOVZJTLpk+lnm+/1sM6879ZvsdxTLxUNPfxSK0nHdpHWblMZStf3yZxf6U9g0pnLUJCnQQM40X4wxaDA5TzuEGogLVAULvBMCr9IHt0iboDrZW/rhz6OuWwL4ybWYtpBISaqtDxWJs1X37q6ALpBoDlvBAaECwJaYSIK51Dhh0CNMfgBdfmDjvYGB47ZAQEaKEKRrAqd7fqKffm52XjTBe5vDURUneSdMQuum6eGjEiw4Bx6Etmfrk8yI/xoqNEkNoxPpyfneqfwcSqjkUFkAH6HT6aoYHNqCs42NbdpWssoT9a1q9Gpayh8rnq/yoA+THPBT/2WeG/GXeYgNq0hm+BVSoYfNBeZeEHIrn/8i035572ob5Ih9Io8XVqCjZ6zg9mm5fybLrCGDaZQOljrQEQ+gRlpUirstESjuM2qxukOnwrzE/7BtZy6cC2R7mFvEJQMOPU443UxrFkotN0GEIPRt5fUHVxbwVthSVt2bqb2gXayI0GgjnbNr7ZyT/s77E6dQbvx8bYD8fTnttCUS8vFLNSiuh5Y5gsuNVGQCZfzf8BRKgtaOiDQ/JwnXTXAeFNeHjSJxdO1iQNDm4vFVAxb3aX4KMdVtLUBtilE4YfWO8ZLZVtmX3tAhufprhoD9H544J5uIcj24Cv788kE9vb/XGYkhEhXouSy6M/Cp96Dzs9kQSb2DMF9OZ0d1OAkyJVQx+Ounz0owk5B/8g2J/42VaD6BJzYoiovXGvFf6EQOAq2R6PKgLOtR+m7GncUtF9RMuNgpPjm6SwiVOMvgPHRFUepKkOg9tMYm0WG+W4WBRtH3/ZB7VXNb4VlqT+C/1z3cTmKFj9AZ2cwx6o1Br/xVUODb5Dr5TNRTB8dmf+fqQwDOKc2q4UCZFtTtdFJqV7T3eM4s/kUJZaxxD3UjqQfJW9H2CMgFN20FWAeIgPLnxkWlXtjVhUPWb/vdkU3ME5LJpt+zJySp0ovoY1jji4F5yAb5y3mSCwNt7xqaYn1QlUQVHftFMQRhz2bvRL4AejA5s9IWzNbebJayFif5A4RhB/vjch0W+3O5PoQtkQmItDYjlhdZS2zK6Qvsj3HpJ9ulhNPnlpQ3+u1pbrE/F4jmmYpNyjxs02+qe7TwrFhpee3TNw251Lb8I/NWXh4koSxTO9UiAFLA+aRrWPoKExQVsLwBKNCwiI50Sx4SqKGyQ6xx/oKIdZEf4RinDKpI7T7IHkSLveDfkKXvD1ZsuxKhAFNe37OJWeep+M3Bth7Ss7upyBwfJdjqPcUwhPbNA9W0Y4WazNBjEVRHa97RnV4ZDWuWM5oPZFylTDt2LibUcRMrd6o79A0oqwCe/vx2RGKH6hky4KlDl59jBrTtXKRh47hDQs6r2Ox/4DvSyDxrxD5kIi6ANHdVUruMd0mUg7zrgRdmwvIuUPFNSzKNzZ3tpa6iXc+iWmFWTQ+o2XoQZWU7FtzlvjtrdIkeuc5MhN+DBvCQMRYBa+3z9jmLm6P0rc1oDakTq5ugmIj6tzoWv+KNljal8iOYO6jqWb1SrMNqdADkCSpapf8KVvEPSlXv3rUROj4Wt5xEejAMeka+DQhdadrqPeTgEAybQaFAhBbhzvMCfkeSUllJ70uidOEbpJdX23Ls6rZdgOnXfgdNutTrl/GIWuY1Sj9IF9ycI1YoRMlq0GBeY0fXa2lYIMce6JsGaYiC7hUXOEPRqpGaeV3GumUhimhVLHQBDzucNpoEKsjbMKUYNBaRZBOAKzCA/OrqceLEThRxwkwL4tuCfWMRaGzBuQWzLgUAHVEgunsIxmj6zOAGlExl15f7MS9JycVJpyh4bv6Q6ieqFRGFhNYZRGZKq7m6OIrt2YhdE18XECznivR3FY8/oMezA+xet4h4ViLhMzFVFtpc4uKaT0UwsB0CIRvlfiEqJ4o9cZKzuNqi8ucYvUoNhx+BxsKaFB0G58SfD5ZevwvXbXwKaWZKhNlpcr24f3BohPwNS+Dzh76AIBmKPYRld5wZcAY98rcoak3+EJ91hyEjrdd3Sk9WNMG4sTufnnN3RLU43MdBElLhnYDOXMKrANM1kuu3IFEPiadcTtSnKX854B6nvvf0vwJpU7seJlZ5WAnb1Ft1FgMnvI0wjSDy42WtNqrNqnFqI3Wz0pQHXqGB5RUdiwua5o2vJyrYZsQzSlAVB8bLf9nvSgwctHw5VV/bJu/13pv06jONjMwJyjdVCQh4Ebsw1gWOHdD1sCRLFJ95i97RF7mv0eJoVO99YE5XkkPUisOnx3QfLDgFWlZKGQMV3VvAvbhzYKYQgCEeTRZgkj7QTURJE00yebTzKodsS0ircgVG+zXgE3XnmtLt948NaO66AcAY4bHEmh3u1zEEAi52oLi9etG9Zc2YT3/X4B46uaMOzy9jZAQw0fuzT2mKqtiCPDAfeGOmOe8bUFdV9luy2NDXorDQloOsP78253hdx4wfIl/9yG4jT0hKXz7zCBU0f7DhqmTdDsYhqbw3vB8qZUdH6sImCdlj66lWYqrCOvTKvPFoh7O0sdMFlbZNmX2oIjJiAZ/CJQ9NtVbiPaHo2mJmRjlIb0JfAmyJxbE3iQCwfjyjNenWSVaivaWodD5/crWvUEssChvJrF6UG3Jx2DJTmOVxvncXYKVbfJ8vsrKDw3uOSmJysckvJRnOVl+vIkT9+r48411wppGMpQ0lP3ch/IT1pSQoO93qyjBiGzPJlUHNjoyv/bVXarZOmy23wlkXMlH8r1n+GC30Hmg3cU00dpPwUi27dmYNRetkqT1cCZuEz7QjzA5XC/K1VhUJZup1wtZ1m3CayO1H/xLK+kcH6bGsuA2fkDX0SIflxpzkTRXL1hkn5LcvfrRR49RwxVxmj54Qa8LuS/7WIAn0Ta5tI6i01evLI/PtJifJY4orfqdBuxZltepxtUnV/uR43zmAQy0ok/qs3AhR3aBviaBphQWx8jTCfZfZfBc8xayZWPApx+YztcT7ArW9hmq1eGIaOi1wGkwAu3Nkc+dPAhLUbhe107vpTp+Arb+vL1wfOubmV6us0ZmXb00llAGvKOAIlRZac9/J2nsHLOEuKZTaZN6WqzkMIvt9EOx3OWaES1GLEXe4YUIi99wl/AjmJyLjycu6/MVWVTM7fwI+HNzFdOtXxlq8ECSti9oAfH7WEhm1LDqBDvWQ5aN2zbFBoqCJzETNLO/hOIKGWQBeUF+iEGj0M+Z1mUcxOyKU7h8xDnsLfZWQXzHwbwCaE/RomFMo/utnUNyTOt/+hs8JMkyOnEYYGWyrgbYa3nr4k5aqrycD1WCRtnrTMYZKyRrCXNi8uvdBkC70bFbHf6sIkHSzoIvdiaKqe8YVsKjePfFUfqHvkzd3BgW9WR+NW0KXOMl4rPgYK9U15KpJRDV3AnjBQzRUCGyWFVh/MeS3rUCCgrKvqpY14c4C6BxR9cvCRmKeTzwF/Elx6yQzDPhwnkWy5Jl4IsITlncIwXSbr0Qw7KPdkM5cQUpkHz2IlnL0tOqNw8qH7n7hCkjpxe34BN/tzYUrCQ6YzOHOoaJwIZfCJ947nYO2qT3FJ6H/NyPyBu77QWDHEfJib6W+MpmdFFrzOlp0wWlxuPzW9AGz8TEsA+c4AFC3aq54Fk1JehhmGlRboyR1Z6uCPvG1jo3nEtHJut6051CWHNyW3eedS+UP3PSJGyEblJ9x8UFLojuqBEkbJhdF22gE0iQKmsn290zkRVz0RGEeCq723Yxo3+rkpF7yDRpB+1wpaVKg7azDKIRg/aOKt8nFSS9TvTo0pE4X6HdzsjNirzpuGojZbUXmW9zLnIznbz96wTm5Audi/21a6lzOEhm58v+t2YOCPTW7BunixpacQFBd6GYFx7kuZn/8JJIR7+10mpSXvjMwKNMzI6BEblYnAK4OrXQSWUsDnz60z9PvvjGMUfy6Il0a95EKE+JwZLp1DQqqLVCmjtMqPsYKaxbMsCvNcZVSgrQKY26XsojcTXEhDmEyKQMeyrs6HZGHEXTFRdPjdTwiNCJ0ld00OQWoyUb7xINsvgZ5vzPRAeO0DR5N9kZ8taoZalEeuhLj18GRbI+61vWFibkVVL0Y9WJO6bxUQcyDeDF98kX5/j6A5Z3QPoByBtkO4rG0eKjw9qnr8Ok/MYqdjOGbAcv85NQtyQxNmECoJAy5/RpsPjqKP0m+13pHkU/OJGeGZp2JoIOpALG14KbjGHQVVHY+Q/ISimBGfEYNdBCJliAMM0Z6il4W1EHZb22Qodr3Qf125cTBlj2cryrtS8GLfWXsZu2nXzoI1YZcxBHJdws3jopcrPqN5SLXBG7CnEwd2fBSq99f9O2vPhT3lm1j4laH9jOhM6eTZqWjjnUVr+gUxBkbEcsLvrxG9pE+IiILF6lmV4GQO0s/06h3qVZRg20QvL4Le9ct71+9J3YRj/aHoNiA8Sit+SLbdUPH2hkRinAbyCYVoivf1j0JCIuofmmk9Qz4ia+uRDhPOgZyiSU4TyP1DGC+LPlvmmEDNS/3SkPmxu2yfTpt1dUL1wos0KHhw1plg/8Fhg4DGR2s3q+hlHpG889gIjNgq7eGKSdyX9mJLG/LOHdigEHCM0bK7luQV6/VP1wRBShrPkKrFOhsV/mxbLTgvYZOczlV+ICtjDA3oJGaZSE4ElHTPH/uDFRO8dNwsxTTWh/su2rXJQwzvkYKdkmGHw9ebRWyjUahFmCjZoRMJiKrEns2V9v9YLOaKQYF24fUEM1JieTxmWfxdNb93t4xMD5LrJAXFFkwMVJ4MpSoSndT9dcNvWeJwWIzhRyJVMSVb2JaGaPYx0RQCRT39NQ6D2HoKW/HMAlNXDFZxrMjaOf/BvYNQkQkZkgn0MpyoI8AH/5bBH9uRR63XaT1sDD4d1qcB6WcWUtgUCN3xyLZCk+dxssQCi+5WDGT0gQIh2tD0+TLlDllFKWIbXYC9g3EnfTiF0suIn6tSjYkQsQvaKtq5hwVf57aR2a82qn4/2VnE6Pmk/LTFQJMWPG1VzgfGUX5DHmVSQEfH2EG5Z2GxdBPIxCoyz6JaDHiQB3jAtKUk7Ti6Qz7V9t8MtRYkgyBcxPKbTvpXHEJiHxVMxQVtt2Lo9axYQo7EZ1EQH0z2xiNEPnQYIKrx7gruKZRNDhzaiDRAWb1DldA7bnUyaLEt7LkTbj3Y3aBW77MgzCWoUlSf69mdtioW8jtzhqGBLXUiDt2JyLw2UwOTGfMgjb1WNBBbQoDZVpbvVkCA16LFytV7Kj2hg3tII5ecENUP0JljJbGOntJrLhC3X6fAvfEnEuESABKfFi5P1hwFmP0XfgopR89vhvThDbuDKTXxtQ6p6fLMc3sKxW9GWICfFhAadX8gNpaC65DH1UIGOK/QuOACPwm5BV0ppRJUhWKdULi8SKicrJd3wNDJeo4X+5/7W0h8SuPfCE2Axs4Y2X9EE8957pjwTDnqJB2SYXMOA29kExYpsZAw+8J5h9/yNCBmswG7X/W0rMamSrmm6XcjXPo2x//H+FiBWZRYHVKFnKJANXvCGy73d1TM5H7GEKdCNRx6fpl5AaxE2XNuDxUryjJeIRGaQGDPNIOTp1lOXUC6cTxVd2cCunCbp0ZLJGsrQ13zXvLv4c29Nby7iIPXAESeiNhNwxiJVN/4jLQ/c6y5FVX1FJ1kAVaoRMZAK1r/Wge/rvQI6iPZ88MlYeEfO9zqGaEu0z9h+qmx8hllNCDo69eia5+OgKo583fwH4/vLp/Y5gYeWDZD3i0oH4sngUh9vqUtVqa/IVAwEaNuLJ33CQtFzbdFW9nVU9DjleD2ijdEzblLCjy87CVvOVLSwiFo29wATdcs3sfBVNP9gmhlUvS2EkXFJU+dnL5xXx87/GXx6uJFTF3/pDUmOqMLqpKbvVZb1B/Y5nh0j+eJ6j8HQmrsf98DsHWE6YLoLrj7Ein/nNFXvvtVQGObHj8+YZLuX+875yCoepC0xtVo9uGnA/ukoFrvzTw0K/X7G287Qu/iK6p+vkdA6dvRsJ7RumSc3yX0E8gGLMOD0Ign2J6miOHFkg+IIvCE7S9uxfw5l9mtDRB3CEwfUGE/HUg1wWL1bPkgqhP2GII4M0SaUdK/hIuP6w1WdfN5jHsI0WqLe2TYDegFyfgnayEP7FGHwYqPNZhov5Tl067tTVbZamAjbwgjENFmJyZ9iH7RYGqsWsxowTKdr8y3nosPt8CJsh7bgGFSsE9nMcoTjpLN3SsroD4LFXasheaaoZmI0VgsmytJvz2Q6TVqAvCEzWFe6ydiGFEEhfQ1FMQ9R+EL4mXZqKn2Jeob2iBSew68kSg0IMAliTOTIeo2U/irzfPuJjT3hYqW9yoHCmqEasJpbFmzm8tPcEPY/ndyBeax1ZovKbVMayZ2jKH0RPZfU1pp+FdozjHNYAE/gSYYkzRwyPlZyrFsjpX0ra8g/R8nPxVe8hi0bRvH9UigXrm9B4T4V/wI1YjZHJ41YRQmfYTpQMaKhcTFShxv2xAqVZ2GX+JWxx/hutNheKfjHU/hJzttHMYBZbjcSFS6Cu6L74LnaAt5f7OeLeDg8MCAnmTS7yQoKkg7Sf+iIAnaz4glA45UgnvZiGpJ8g+4lBG/ZZgXI8ETBOccJH0UuvdxWdhLE+XvN2gLIVS15u8Ahb6bJ8n8CAKnnB1hpt3TX2d3iaUZORToeB+3acdr7t25ozvfaNEvdxZVszOpOwlNUBRyz4X0N4ArkSm+meDfA4SXNO5iXLX9pN3KwJnrx16wGYI9yx5PphWtI2vZpa7uKB2kl2O2aAkN4ITiiPfvjyAnROZOgS3ksP5I2n6tF3av6FHSl37BBLsR57Z6Sh2ndM9ON0uGZAmyzX57yYSmAK4rURPDBdxQu9RFl1sslBwDOe2v8du5Nc0Ct25P1GnNgneLGUeiUtRnWTD/P0U1RqibeD8d5G5iEoVZyeFACKzqo+ePFhMOG2+E1YjHlNX2HhBML9b90yFNpDm1LZj0bbV4spDn9oL7ipiJERbtLSQy3sCB0S4Tu+5i3lr58ORFUWi1ToNdUZq2bBx/IE9ZfinN6kpip5QOjk8+VJ+ZrRS7S6sCr4zfpMU6XJjzz0wVq8XD9PbmbZGyj0TrOsr4tKNnF7Tspqfj65BdLg9qDc1wspvaZvb6RFO6BHlPAdLcCvcgwa26ctMgyP0zO03phLmlbl0fVDe+AjcpSmWJFLxXIJ+UV5jrbZQQBMcMuqFJFb7wCF+4wAT4Q7rBnDWsdjHkgoL9Fc8c3QlYF5ZUcIRLZmq8InB5SC11KbGh5Cp3PqTwzne4SEn3JoiHV//38RJFGUyGhf8n2uIfd2h6TkZOXFhEkZ1ZhYL2aSPjoCzLyaEGUFz17RLyqptrVI1hCO+8N7KZ9nxNW+JYgpwVO2LGY30ch3QX9tsRR1AYLIIo1tvmqOBbNiLL1Bm1+ieO/aGyputXLsDZhgaNihZDJVRKWaWpGh8bbktE+1hBUp34lQGk86y8vNUYikqzPcgGFYjS3zsWvunmHgF+yPy+mz1lbHh50XQUZTwAwmXVXRzYVulRdf0IsiV6pbxvyNv/DrZdPW4syViT59gnPuMULuZCQgArwQCvvbgLffPcwxVJcQlDmr3DZdV73FV0FX1JY2tDfb1GrUqw1+Z8wOqpGnFWQTuajox4eCXXWmKppJ8izwlmuPPq1aTqShCOmJyGGPKvnf7lDY4QPCRjqTq1Vu1IEcMqj0v6QfXcjuzjvCWGnswlz4C/bu3Yn7N3eHfFVp2I5X7UHHFr2ysuXYXJCChp3Rgnw5lZFWhPZDtTpMy4kHPfhaeopdEhAib2AtdlqB+Z/0Tt0RvvZ3EFkIlr3ySMbT1IlRIYoUOnhl/eav9rrf6AI80DSZMm/8CSO2fr10tg5vM5xoG83fB0v2RRIPc7culBr1rn4Rwhm++PLcBBMMtQyDYaCaRN4CpgvbMsyYE+TcprYHhqIgq3t5yEmt7uLnQPiqwePcfqCje+731Kj1xvI+zpvcrOFTiQToPhFL2Kjku/wOw+xPmmhmkI9128BJEI813ejOp7EjX7myTHzxlZY5kcVRbxEdvI+2bhCaZVKMPx4titnF/HehbFDqR4jGbemEmzp9VdQNB9O93U0t6bhZc4jumz+tB/PwX23nyhAEufJnoCKl1gVWv8WVOvhU/FEWw1jMAP282no35rt4h5LCP07/+sf75KaYhcpMbAEj2xbLhOr4DEDf9zGak51u5uVXhBmF0wrkNT2vuYHfZjlT7o8LpyM/vmZ2Q+I7VAKdBALprRj0tF5INz17e67R7MLlrCKIF9ta3vIlM/CJqeXkNh+tlmcnP6qRWC0VuIjIbv1Qv/rrtRrAluLlXesmYeKiE7/KXrWsgikJ48oVB26FpfdG3gXbf7JQTR7tED5y2vu9qZdQ9Wdpu3KHVbgg+GA6AZg0fylfv8YaZHy6tuk05ldzLiCrX4e2PNIfeLwVKW+0lOTByCWsgOcOJiQeiew74cHY5qu0ovA9unBzRlT0QOeAc3vBcyJNH5/SWBTR/8LUTfKeb+Dsy6EPRiXIeYGOPq/+PhQj/7dF0XcBnWn4qjsvTquDUbQK2VhpjgJIMCHI9V3p4hW1lhudQeQN8iC+hqtAopBKtuwkx7Ed/MMqtlAg/kv3IHBfqJqqZiu/Kmk3AyhaKb8XUrUzJ9dbMBiATVjcZV7xnjMz5falEe4eVy7xGQjdFx/jynCtws1z60hLfOy8I2CkbYfO3cjLoRvyU3nxst3KNd9jQiZMWVjeFqJ6TkKAS6Ir5ykRbgG+bsDBqXtz8ERVbqRG8Xp5YZyGDIr5TZSki0Sfe1UW7Qmqw+JoUeEfthJ8AiNSOpAU1FAyYSo7tOTpg1izo8LIxEikC1/tocbi4qCwsoFJgaGhqoJz5eDDGvJa2wTjjtmf2O7CbQIxE2lLLmmMjx7dIIk4/4m/3vou3/3SPJAm4imoIOEDc/cVYF99f37mAspzFSbN1dCqPfFmbP7DuQW/KD8ooMx/ID4/LOzk2lgumHh4Ajo5kUb69t9Rcsm3z6/g6MigdicJYpZOBr4iKSeexeb/71847SfuY6Cu6cn2uEpdSPZRW06kW8JRuARSjfoClpH4gLTbfiTCNgmDqU+S44wRKvF+YyXlGwsE7SCBVnxQuDaeyO8x+RAkKCQzblAi8Eux5r2I1QDvcMA4gPxbyO1WNeORSF/EcAKI2+cHlQUHFNpfi79lU//2n0MKeg3RBbph/9xY95lfNtEj7UBtVS7P7UgGN79jVnv4GZhrCclXz1KEGF2MjaVAPhVPrFfS8g8LTXw1Y1GDDv9z4aR3Sb76nHJspZiUHdd4vdqaD9kbiFJLEzcBjWp/ByuAuOePg09c7ctP1OxoE9JzC/FdI9TCrmtGuuFWmcHpa4vrmYlB7sO861QPqSoiTKuKzGNMlemKu17k5umKT7qsRw+tNmtWFsHFek6w6RaFDaDiYWfSc6aA6eEOqUJL2ImAISi6wGM3trDc9XeAaDrYqt5WW8nfbOjHVVEoof2MOB78sdAOMQGZpSniETtcm3zqg3m9RvWYrJV2DGnKb750wyUa8izwABNwdWJ5zJFaMi8w+Dq7XxJ3zNLDlfiTIPhzFAg3hSpLX+jviyLEMhsZmrGUCRq/EeqvX0XjA2/gpEmTRORUgg3oKHyCcXVnSo5iyq614r4O20qe9fxTYDDKohbAE7EckyaBqMLZiiZCwrmIqWi/Oi1sRti/vf7LipOG9YDrOXGJWJ0VKBhJ9375DsqU2x+VFoWlTviXr4mG+tAexghSA7qUn8m0WYu1Qzzmo72jsOZrDOp1/fiiU9kx9zCx1MtLB0E//53Rl6bHjok2rbOkzPJT0grWC5WkVqPlbwXufA7N/Mcorq/oBi9StB9IGhqjmh9KcKdOPpwTkojWqnCpS2ZDWqGiWBwoegPSQDV3HeNKjvS8BMjI/9yzHZpZk2RBtaFlUohhUgHf1QrXf/OFSb9B4IzKTh8dKc3+n+siWnUJL30IwewK/pmYL0ZGn+CX2jOjkx019NNPoB8T4S5kNKYym75cwKW5AvU74M71NwRk1OffCkd+rznWuAhgjs5fkzu1IptQmFHS/y53jRaMC1FamrhHzNRbSgrDi7PUxNrZpThUzH3my3QjozcmbzxKy8RN8rK5msof+bg3W5Sv7qYMxQf2jLdbUMwMAa1Wdx/tdLDFuQrK+eTgqg7ZCqrNG3DqNBk2aQjCfRYZhFdeTx5hVEyFnTxfvzH6gmbmXqFss60odBpA7uDM35nd9E9SJsTT6hmWT62tIb+Z/PAWJJWAMAEzuKg9FdjoSdsYPS+G6Ks7N5D0ONSwxu0t9CRfHBfUT9fTA3Jo2vVzhuK8Ki5kJsAqFZKijIfEXi/66xk+t2ng7q+wYiPUc/zIf16RJwSmbmzFYsVh9U2MwjmmyeaaYC6ijr0CQ6Lir3rTn2+nvNJxi9qS2fra3FOyg6UNAXMLfj881TuBfSf8nxdyHfABAyNAwjfi9EkyKHpCyg3e2wiAitfnVoNh4NCYuqMI/Y3McbtQ1B6xb6BOyq7UKJkqlZEFfLAURa1WOicNBZluNkMdjXqJNBXC0sBfxaEaNn8u4zRnWDR4JYWSkxqSeprqYoDCRW3Oe7AwlNOMG+pnFBHRvwfC7wlp9xS0yC51gBbUyZVx6+8QPrTHrXyYIglu7ZuNqofg0Z9gMdbyxO8hZ0Fx+VWEPWvXYNlNIOpeGlBbje9A5AOWwKS6vgb58vvutheZ2cT/uMjOfQB/qg99KUkAhXjWZic2ucFpPh1DgSN6scS/CydTg9TPL5A8F9rhAU066eXp21Xjf7yzkZf5+uCtVZOSxV0vewd7OjUqm9pXsKxMBXTkzmsmCIAC/RWWC4HUZawrAbyF9sRzUCOSLuaKgnwTlZjxzOQnVpahPauwHIQpWr1GOkvpQ40NhB4PdrZoKv+GESH6Pls61Mlf9RYEz0yrxu1BxDLE6rAVHTFggN0uZNqcVTIPpoT7QnXMRzFZ185ABuF/DWFXV+ChKG6DogCYTPm0gpsFO3V7WR1gdsRFFtPBMZX9ypTMDhrvRz0zzSXoJAJGwLvdo5t+IeTbxNEmt7GpDKJlOlKhn3/+x811g2gCDvnhULtpXb3K7FvEw8brBzAAeR04LmNY+Yi5DkpLxrIBaCkPprcN0BQPq2TDYFXM6WKK4tCWr8CmWpXPxPMJNfDVyxeAMSTGamHqpDxf5sTfJFXV3AAQrI78pLTvad0WkQuuw2RBOz+zUlrqJYsLSwiS59Nt3sJioI6ClzLeGFlP3qjQ9LOeO0xzQ1eGLU36MIjpMB0+wOFKP7TknZnS6LOGfHSAjfW7cALIAltt2b49L3X/j9IDRoO3VhIu6A+8vVs0Y5f0b0pjQCEq+OOopUOkIXQNwqnEtKQfC+AKZ1hAJfXU7R6c3O49ZDbmWYHTj/I2Ql0H5oJn9RLyDg1GhmAlNcWH/cmPCVjhk1oND/qzWdJ/zkyO3r0n5FqhmO66pf7D9W6edIupjHSdS4kd/Kn8BmmRLpIEHEhXP0b6Xdw0Zt00kxPQ3WqjrQsvDhT+ZdAjAgMVEcBznPt0YzhTBFYwrEBvYzg0ly9caZ26XfrGBckZE8SHCGejc4sMvA7gY4utl0UQfz8uId1F4BePdNA73Hh6Kp7e0B9zhQuxk3XyX++d2k3TjgZkn7tEqeUR3bOCd9n+juFVS7bpHRSBZfAou/5duzo7Fu9XP/7pfuB0XXjSA5yOrcAetqNFoTKV7SqRlI8Ogbt8bvnXfqdzK0X6NnN8k0C8ascFzgmyh7wwr93Tq2JIDeOwlBOtOddt6E40XdPbd+JL7lsOiAp3LHq5X3KVe6IHTjcOhoJn5ILIAFe7BtyHIBYjAuw/5T8asasdGdF3FlmMmyS002EBofRuU3N/H/LTSzbTukBx5l9LnJwfqM+nkBfpHZSVDPyhVdtWxWW1puvct5FMQix8SUUvsVsHbeB8G0CdiAiiiQ70t84rpZGmzstWwGE3WFyk3jr/NTHZY/yzRrXIbF69bKWfkH9SFrpIBJ4ifOTtqtby0L93aFLHPyFazc7yqWpXX5GjH8e9ISFIe6CVgNF/ySod8WqQXYUCUVHNX0vn1wPRY9hEVxxOnRJ/OJFFWjcPWzah7Z6Y+XkLGDTCxSFs3qsfFdCQEbA+kJhtMAXLqSpUyitV8SItjTGykNynyWH2Yl4cWH67PO66LtTBhIMBGEX5fXLErnGmZX+Gcz/shEM3YKWcNGymOhiBFui4zTa0MZ6u4WACMYY7H+0aa/lZhdaaum+xYJTED0p9N1vIraqj8PZoRcgYwt6CYFf0U9ZqW5fqIVHfnEqwutx/CY6McoAGMSzMsDas93GV4qeziVc0oMyJGVIiax4DdyOMFLVmjYqAKPAfpA8GhZd6J8ThdMIHRz9jKImqGOcHpRJ4JhsQxLpZnPJJeyRu2+Hd3SD4DZ7g2DWGkUduCrYO/URbeunaFYobXPMI+yx82856TeIx/yAR2Q/zaVzQ0dlQqDvuBE5s1fHqfGCcNIo1sVwoi3NNEaXHW7MTgE7fgzX+9oGatguDRMEt2XPVkV3CJSrOZSWCC6uM5vOQfPkoSomzFYkjetSRjH1ZMu9M8XbWBp/OIKZFHKmjN3wcaVfSwK2Y02MuBEHOnCkuc7xNAG9s06+xOImNgClRTy9doZK9MSuk+QW5QC9P2si7J2h7SPn6ucg8sgsYLhIqXlHAmBfTYxNWWwsTb3WayII91K3YimFtFI7co7sTvA7fI2RMshWJHvfotqQZILTRoo9JKwW+EDdpkH/iwy0bSkdHWutsEU1bBe0KpUqdRWdcrAwGNRrth6iN0V86Sf5MKzGpOQVC+wx+VAeKw3pKjjuV7szWux33Ga72DWrLTi76l1yo1MxN59IRRiDQVmBgxgiBVp6Ieh2hzb93/HC9Z0n8MsPVWVbuAQEct5vs4Q8Zk0VFUrFOAUlZxecDHpCLr7YxtMaLvSB2o/RDrUNFt+eywnz344v30rFtjOrsTxs+HTQUtajpu90KqqDcHbx9MxQfjCJ2AOKQjsoC+AqnFuX7dehflIveewlbOVUdwoL+GV74V1FiqRw5He9wbSIE5tMrWfdN0FQhStmzEcEhup1GL5/A7JUaRUFuO91blsO9Wtht3vtcyBZY1qobILgkzQip3Mt8lbmAXNLLcufuZqrOq81PdS3NAhSQRpMaEV6uiWWQo9q8wyho1+htgQUk+YBFXOIDJVB3vWegQSt28fTbaNWHhpR1XVaG8N5H6wYNkONg94rp1TOGC8TQbaeBSGNXdL32rny/TRGgJ6cqs4iqVR2tXdi6QDZB9cer5lp7nW7Y2HDupk5THe37IsWEDapoYnIY0dUp02INILN49XCqFHlTVhbiXgmK17eKH9vKoxI7SiPRW+mxZcJlrjAkajiB6pPoFpPAUcI2nMQYr6Rs9OJPNyynhTT4GFHmk5u4BITeV4+Mnh3iDq1pohehW88d1arRYOAbc4u6/nj8oDZno9pEUnE7hqn9cLmRbi6ZTVgoC71jX3pjwU+J93MTiVUuIiFnTp12GG+hTA6DW1PAmdeDraVG8szWPNYlGTXqcPuTJMbg/blUoqBg+jve1RfEVXWCiMt6A4MYRl3u0E8gz60Dq6OG7WyIEqWCUUaA9cTyZVrH6keQyk5SJiycxjwuhNocTS46c2tMkwSjhFGPPhV7Vv3B/0dKZ3kUp7VYxZdGDWO6tPqwvV/H6JZQCJubCjKP6iuX3uMIAFOMRP5IZ4zZKEh1IkNeRdFyYw50gTeQstbGY3GOj82Gmo9i6Kw6hrRozPADeWlWovbi6bQazllCVHYoX00mBV4hvT/95i2OscsjD79ZyJdN3YgXt0PVNVxFKBCvciwjniVtc+jmRx2pRBvXrMjcRgIDFmwsFOvJhH4HwtJVkQ+M5ZEM52ihZ/ek0qdFd6gjgbbTm0lsyR8WWcZ1m3GapBTY1ZVFd8CDn9vvShSvhxdlvym7ZzHX4D3jgASKlhi6R1p3Wny+2Iuh0ftM4upQpYRR92uYE4DdNW7aRA2CwFLQRgIbyB0/1U+Lpabx8gI4xkrdYE+sNNPKAVei8WJdLmmi56Sa6XUkK7A+RjNEgYG12AJ7CnjzC9YC5elR9YyLZ2gG6JiORFE3ufMmXdDk+Z+cOoLD1eQuYbaFrtWh1W3QtSKU3qNxrZ3Tqb2JOdSzPIIvj414NMscC6S88ByfcTIrT0DpDuYh78MIJxcHh960tTF9hU67dzpHkqW5rwqk2Fdn5FMzPjeelCZioHjcUGPq7NaIf1TG9YbevrX2gLtGHioVrGJzOKKccbqU88GK4IxV0Cg+kU11RS41WWYDUYMis7gase2Iz8y7Q1pBkceyea/EqoaYwNIEmnBm7NP1UJX0yZKQs1wOw6d9uZiMDPrxG9rRUY7DE7sGOnlqQhIzkGBfxNihawqwadfAK6jxw94zHPiH5KyIcawCdNRJEOPmGfFdC9bZo6FJgh1TJPZYU3kH2q/TEqHSpQElaaWGbb/t5HRhJzNz+wQS4X9ibeUa9heaYAlGWMjIROdI2QwUZmdOwUTtFALYaHO5uyU+CntV8w9Y1f/k7ZVtGbgJjw+r4FSK8HVd4536Q80Opu/cl6TvfUvFpI5KLQOmWPg7ER40KizfZapfjmSTyIgvKBXICK/snIGa4mEshwdCOFff43TuKf+cIsfFhS4WuxrJBlAmM1dd4P34zee/FUnyewHX3a718Ai+0B7kF6qII5f8Ke6Aj4c4O9R6lUa4vHCiJkC4hb/+UMQnLOLReJCIuZzKyue/h4hfw+kJt/Cper18VLPuIsO8OzOdCURCLE60cCzoyQ6QA74TM0+aEU8R3d4q4r1osoRk53fkG1Lv50YVnHRv1PVmx2IG5WkExvQekDby8ojlqI/m2Kts+jIxQNaaQzndXa/giZwyKhCheUtlhCWXRyzMGwqZpZS0Cd1EyL/mniU4MCzJGsPb8Y6d7qL+zFYlEjipBa0qwG07nF2T50PDyjQV3gKSaXc/uiOZt3BkV4kFHhsvttieaTV6cO//RlwMsg2Nod+8xfyjmxXlhFXX7G2+RNqsyEJZpM/ic3LGr2ttPv1PHip7Df+Hq8agpgjVJu04DLFqa3MIMspDzezWc9P8YncGjgsddz4catHgewCzWtgbJipfdhqH/pYURo7BPHpqN6RtSLNXAT99VzjmZQkO+nhj6ssuBNmcrkvgSHfDabrm/WmBMMDuRgxJ7vhH6YglOoxu111vIO2N4w3THFntPzf7hlYMIW84CbCTrHHBv9bgj7ly0wrHum6iIPM/Bv/yGuZjXRA9atw5r/LihAPynM8ixhiBP0MnjMQS7hqrTpKxSwaG00FKUyFpA6VjGm7GCRbzAxdcIvQ9uV/f09TK4JfMsjmhRaw/qvlKaM3AKZgEx5gKS9PpOj7ztoKdtT5nWWrPAyDU61wqu019nNAbZ+AAt0gwknuQn/cstrNDTQ//L18vYnNjZnJhbWU"></div><input type="hidden" name="bgresponse" value="js_disabled" id="bgresponse" style="display:none"><script nonce="c6XQoK_6ljSIPUPPhVJTog">(function(){'use strict';var d=function(a){var b=0;return function(){return b<a.length?{done:!1,value:a[b++]}:{done:!0}}},f=function(){var a=document.querySelectorAll('div[data-button-type="multipleChoiceIdentifier"]'),b=typeof Symbol!="undefined"&&Symbol.iterator&&a[Symbol.iterator];if(b)return b.call(a);if(typeof a.length=="number")return{next:d(a)};throw Error(String(a)+" is not an iterable or ArrayLike");};/*

 Copyright The Closure Library Authors.
 SPDX-License-Identifier: Apache-2.0
*/
var l=function(){this.i=new window.botguard.bg(k,function(){});this.h=this.g=null;this.i&&window.addEventListener("load",this.j.bind(this))};l.prototype.j=function(){var a=this;this.g=document.getElementById("hiddenMultipleChoiceIdentifier");this.h=function(){a.i.invoke(a.l)};this.g?m(this):document.addEventListener("submit",this.h.bind(this))};l.prototype.l=function(a){var b=document.getElementById("bgresponse");b&&(b.value=a)};
var m=function(a){for(var b=function(e){a.g&&(a.g.value=e);a.h()},q=function(e,p){p.keyCode===13&&(a.g&&(a.g.value=e),a.h())},g=f(),c=g.next();!c.done;c=g.next()){c=c.value.getElementsByTagName("button")[0];var h=c.value;c.addEventListener("click",b.bind(a,h));c.addEventListener("keydown",q.bind(a,h))}},n=document.getElementById("program");if(n){var k=n.getAttribute("program-data");k&&new l};}).call(this);
</script></span><span jsname="ZVfTqd"></span><c-wiz jsshadow jsdata="deferred-i3" jsmodel="hc6Ubd" c-wiz><script nonce="c6XQoK_6ljSIPUPPhVJTog">(function(){'use strict';var aa=function(a){var b=0;return function(){return b<a.length?{done:!1,value:a[b++]}:{done:!0}}},n=typeof Object.defineProperties=="function"?Object.defineProperty:function(a,b,c){if(a==Array.prototype||a==Object.prototype)return a;a[b]=c.value;return a},ba=function(a){a=["object"==typeof globalThis&&globalThis,a,"object"==typeof window&&window,"object"==typeof self&&self,"object"==typeof global&&global];for(var b=0;b<a.length;++b){var c=a[b];if(c&&c.Math==Math)return c}throw Error("Cannot find global object");
},ca=ba(this),p=function(a,b){if(b)a:{var c=ca;a=a.split(".");for(var d=0;d<a.length-1;d++){var e=a[d];if(!(e in c))break a;c=c[e]}a=a[a.length-1];d=c[a];b=b(d);b!=d&&b!=null&&n(c,a,{configurable:!0,writable:!0,value:b})}};
p("Symbol",function(a){if(a)return a;var b=function(f,k){this.g=f;n(this,"description",{configurable:!0,writable:!0,value:k})};b.prototype.toString=function(){return this.g};var c="jscomp_symbol_"+(Math.random()*1E9>>>0)+"_",d=0,e=function(f){if(this instanceof e)throw new TypeError("Symbol is not a constructor");return new b(c+(f||"")+"_"+d++,f)};return e});
p("Symbol.iterator",function(a){if(a)return a;a=Symbol("Symbol.iterator");for(var b="Array Int8Array Uint8Array Uint8ClampedArray Int16Array Uint16Array Int32Array Uint32Array Float32Array Float64Array".split(" "),c=0;c<b.length;c++){var d=ca[b[c]];typeof d==="function"&&typeof d.prototype[a]!="function"&&n(d.prototype,a,{configurable:!0,writable:!0,value:function(){return da(aa(this))}})}return a});
var da=function(a){a={next:a};a[Symbol.iterator]=function(){return this};return a},q=function(a){var b=typeof Symbol!="undefined"&&Symbol.iterator&&a[Symbol.iterator];if(b)return b.call(a);if(typeof a.length=="number")return{next:aa(a)};throw Error(String(a)+" is not an iterable or ArrayLike");},r=function(a,b){return Object.prototype.hasOwnProperty.call(a,b)};p("Symbol.dispose",function(a){return a?a:Symbol("Symbol.dispose")});
p("WeakMap",function(a){function b(){}function c(h){var l=typeof h;return l==="object"&&h!==null||l==="function"}function d(h){if(!r(h,f)){var l=new b;n(h,f,{value:l})}}function e(h){var l=Object[h];l&&(Object[h]=function(m){if(m instanceof b)return m;Object.isExtensible(m)&&d(m);return l(m)})}if(function(){if(!a||!Object.seal)return!1;try{var h=Object.seal({}),l=Object.seal({}),m=new a([[h,2],[l,3]]);if(m.get(h)!=2||m.get(l)!=3)return!1;m.delete(h);m.set(l,4);return!m.has(h)&&m.get(l)==4}catch(B){return!1}}())return a;
var f="$jscomp_hidden_"+Math.random();e("freeze");e("preventExtensions");e("seal");var k=0,g=function(h){this.g=(k+=Math.random()+1).toString();if(h){h=q(h);for(var l;!(l=h.next()).done;)l=l.value,this.set(l[0],l[1])}};g.prototype.set=function(h,l){if(!c(h))throw Error("Invalid WeakMap key");d(h);if(!r(h,f))throw Error("WeakMap key fail: "+h);h[f][this.g]=l;return this};g.prototype.get=function(h){return c(h)&&r(h,f)?h[f][this.g]:void 0};g.prototype.has=function(h){return c(h)&&r(h,f)&&r(h[f],this.g)};
g.prototype.delete=function(h){return c(h)&&r(h,f)&&r(h[f],this.g)?delete h[f][this.g]:!1};return g});
p("Map",function(a){if(function(){if(!a||typeof a!="function"||!a.prototype.entries||typeof Object.seal!="function")return!1;try{var g=Object.seal({x:4}),h=new a(q([[g,"s"]]));if(h.get(g)!="s"||h.size!=1||h.get({x:4})||h.set({x:4},"t")!=h||h.size!=2)return!1;var l=h.entries(),m=l.next();if(m.done||m.value[0]!=g||m.value[1]!="s")return!1;m=l.next();return m.done||m.value[0].x!=4||m.value[1]!="t"||!l.next().done?!1:!0}catch(B){return!1}}())return a;var b=new WeakMap,c=function(g){this[0]={};this[1]=
f();this.size=0;if(g){g=q(g);for(var h;!(h=g.next()).done;)h=h.value,this.set(h[0],h[1])}};c.prototype.set=function(g,h){g=g===0?0:g;var l=d(this,g);l.list||(l.list=this[0][l.id]=[]);l.m?l.m.value=h:(l.m={next:this[1],v:this[1].v,head:this[1],key:g,value:h},l.list.push(l.m),this[1].v.next=l.m,this[1].v=l.m,this.size++);return this};c.prototype.delete=function(g){g=d(this,g);return g.m&&g.list?(g.list.splice(g.index,1),g.list.length||delete this[0][g.id],g.m.v.next=g.m.next,g.m.next.v=g.m.v,g.m.head=
null,this.size--,!0):!1};c.prototype.clear=function(){this[0]={};this[1]=this[1].v=f();this.size=0};c.prototype.has=function(g){return!!d(this,g).m};c.prototype.get=function(g){return(g=d(this,g).m)&&g.value};c.prototype.entries=function(){return e(this,function(g){return[g.key,g.value]})};c.prototype.keys=function(){return e(this,function(g){return g.key})};c.prototype.values=function(){return e(this,function(g){return g.value})};c.prototype.forEach=function(g,h){for(var l=this.entries(),m;!(m=l.next()).done;)m=
m.value,g.call(h,m[1],m[0],this)};c.prototype[Symbol.iterator]=c.prototype.entries;var d=function(g,h){var l=h&&typeof h;l=="object"||l=="function"?b.has(h)?l=b.get(h):(l=""+ ++k,b.set(h,l)):l="p_"+h;var m=g[0][l];if(m&&r(g[0],l))for(g=0;g<m.length;g++){var B=m[g];if(h!==h&&B.key!==B.key||h===B.key)return{id:l,list:m,index:g,m:B}}return{id:l,list:m,index:-1,m:void 0}},e=function(g,h){var l=g[1];return da(function(){if(l){for(;l.head!=g[1];)l=l.v;for(;l.next!=l.head;)return l=l.next,{done:!1,value:h(l)};
l=null}return{done:!0,value:void 0}})},f=function(){var g={};return g.v=g.next=g.head=g},k=0;return c});var ea=function(a,b){a instanceof String&&(a+="");var c=0,d=!1,e={next:function(){if(!d&&c<a.length){var f=c++;return{value:b(f,a[f]),done:!1}}d=!0;return{done:!0,value:void 0}}};e[Symbol.iterator]=function(){return e};return e};p("Array.prototype.entries",function(a){return a?a:function(){return ea(this,function(b,c){return[b,c]})}});
p("Array.prototype.keys",function(a){return a?a:function(){return ea(this,function(b){return b})}});p("Array.prototype.values",function(a){return a?a:function(){return ea(this,function(b,c){return c})}});p("Array.prototype.find",function(a){return a?a:function(b,c){a:{var d=this;d instanceof String&&(d=String(d));for(var e=d.length,f=0;f<e;f++){var k=d[f];if(b.call(c,k,f,d)){b=k;break a}}b=void 0}return b}});
p("Array.from",function(a){return a?a:function(b,c,d){c=c!=null?c:function(g){return g};var e=[],f=typeof Symbol!="undefined"&&Symbol.iterator&&b[Symbol.iterator];if(typeof f=="function"){b=f.call(b);for(var k=0;!(f=b.next()).done;)e.push(c.call(d,f.value,k++))}else for(f=b.length,k=0;k<f;k++)e.push(c.call(d,b[k],k));return e}});/*

 Copyright The Closure Library Authors.
 SPDX-License-Identifier: Apache-2.0
*/
var fa=fa||{},t=this||self,u=function(a){var b=typeof a;return b=="object"&&a!=null||b=="function"},ha=function(a,b,c){return a.call.apply(a.bind,arguments)},ia=function(a,b,c){if(!a)throw Error();if(arguments.length>2){var d=Array.prototype.slice.call(arguments,2);return function(){var e=Array.prototype.slice.call(arguments);Array.prototype.unshift.apply(e,d);return a.apply(b,e)}}return function(){return a.apply(b,arguments)}},v=function(a,b,c){v=Function.prototype.bind&&Function.prototype.bind.toString().indexOf("native code")!=
-1?ha:ia;return v.apply(null,arguments)},w=function(a,b){function c(){}c.prototype=b.prototype;a.P=b.prototype;a.prototype=new c;a.prototype.constructor=a;a.fa=function(d,e,f){for(var k=Array(arguments.length-2),g=2;g<arguments.length;g++)k[g-2]=arguments[g];return b.prototype[e].apply(d,k)}};var ja=String.prototype.trim?function(a){return a.trim()}:function(a){return/^[\s\xa0]*([\s\S]*?)[\s\xa0]*$/.exec(a)[1]};/*

 Copyright Google LLC
 SPDX-License-Identifier: Apache-2.0
*/
var ka={};var x=function(a){if(ka!==ka)throw Error("Bad secret");this.g=a};x.prototype.toString=function(){return this.g};new x("about:blank");new x("about:invalid#zClosurez");var la=/^\s*(?!javascript:)(?:[\w+.-]+:|[^:/?#]*(?:[/?#]|$))/i,ma=[],na=function(){};oa(function(a){console.warn("A URL with content '"+a+"' was sanitized away.")});function oa(a){ma.indexOf(a)===-1&&ma.push(a);na=function(b){ma.forEach(function(c){c(b)})}};function y(a,b){if(Error.captureStackTrace)Error.captureStackTrace(this,y);else{var c=Error().stack;c&&(this.stack=c)}a&&(this.message=String(a));b!==void 0&&(this.cause=b)}w(y,Error);y.prototype.name="CustomError";function z(a,b){a=a.split("%s");for(var c="",d=a.length-1,e=0;e<d;e++)c+=a[e]+(e<b.length?b[e]:"%s");y.call(this,c+a[d])}w(z,y);z.prototype.name="AssertionError";function pa(a,b,c,d){var e="Assertion failed";if(c){e+=": "+c;var f=d}else a&&(e+=": "+a,f=b);throw new z(""+e,f||[]);}
var A=function(a,b,c){a||pa("",null,b,Array.prototype.slice.call(arguments,2))},qa=function(a,b){throw new z("Failure"+(a?": "+a:""),Array.prototype.slice.call(arguments,1));},C=function(a,b,c){if(typeof a!=="number"){var d=typeof a;pa("Expected number but got %s: %s.",[d!="object"?d:a?Array.isArray(a)?"array":d:"null",a],b,Array.prototype.slice.call(arguments,2))}return a};var ra=Array.prototype.indexOf?function(a,b){A(a.length!=null);return Array.prototype.indexOf.call(a,b,void 0)}:function(a,b){if(typeof a==="string")return typeof b!=="string"||b.length!=1?-1:a.indexOf(b,0);for(var c=0;c<a.length;c++)if(c in a&&a[c]===b)return c;return-1};function sa(a,b){b=ra(a,b);var c;if(c=b>=0)A(a.length!=null),Array.prototype.splice.call(a,b,1);return c};var D=function(a,b){this.name=a;this.value=b};D.prototype.toString=function(){return this.name};
var ta=new D("OFF",Infinity),ua=new D("SEVERE",1E3),va=new D("CONFIG",700),wa=new D("FINE",500),xa=function(){},ya,za=function(){},Aa=function(a,b){this.g=null;this.l=[];this.h=(b===void 0?null:b)||null;this.j=[];this.o={g:function(){return a}}},Ba=function(a){if(a.g)return a.g;if(a.h)return Ba(a.h);qa("Root logger has no level set.");return ta},Ca=function(a,b){for(;a;)a.l.forEach(function(c){c(b)}),a=a.h},Da=function(){this.entries={};var a=new Aa("");a.g=va;this.entries[""]=a},Ea,E=function(a,
b){var c=a.entries[b];if(c)return c;c=E(a,b.slice(0,Math.max(b.lastIndexOf("."),0)));var d=new Aa(b,c);a.entries[b]=d;c.j.push(d);return d},Fa=function(){Ea||(Ea=new Da);return Ea},Ga=function(a,b,c){var d;if(d=a)if(d=a&&b)b=b.value,d=a?Ba(E(Fa(),a.g())):ta,d=b>=d.value;d&&(a=E(Fa(),a.g()),typeof c==="function"&&c(),ya||(ya=new xa),c=new za,Ca(a,c))},F=function(a,b){a&&Ga(a,wa,b)};var G=function(){this.g=(typeof document=="undefined"?null:document)||{cookie:""}};
G.prototype.set=function(a,b,c){var d=!1;if(typeof c==="object"){var e=c.ha;d=c.ia||!1;var f=c.domain||void 0;var k=c.path||void 0;var g=c.ga}if(/[;=\s]/.test(a))throw Error('Invalid cookie name "'+a+'"');if(/[;\r\n]/.test(b))throw Error('Invalid cookie value "'+b+'"');g===void 0&&(g=-1);this.g.cookie=a+"="+b+(f?";domain="+f:"")+(k?";path="+k:"")+(g<0?"":g==0?";expires="+(new Date(1970,1,1)).toUTCString():";expires="+(new Date(Date.now()+g*1E3)).toUTCString())+(d?";secure":"")+(e!=null?";samesite="+
e:"")};G.prototype.get=function(a,b){for(var c=a+"=",d=(this.g.cookie||"").split(";"),e=0,f;e<d.length;e++){f=ja(d[e]);if(f.lastIndexOf(c,0)==0)return f.slice(c.length);if(f==a)return""}return b};G.prototype.o=function(){for(var a=(this.g.cookie||"").split(";"),b=[],c=[],d,e,f=0;f<a.length;f++)e=ja(a[f]),d=e.indexOf("="),d==-1?(b.push(""),c.push(e)):(b.push(e.substring(0,d)),c.push(e.substring(d+1)));return c};var Ha=new G;var Ia=typeof AsyncContext!=="undefined"&&typeof AsyncContext.Snapshot==="function"?function(a){return a&&AsyncContext.Snapshot.wrap(a)}:function(a){return a};var H=function(){this.I=this.I;this.g=this.g};H.prototype.I=!1;H.prototype.dispose=function(){this.I||(this.I=!0,this.H())};H.prototype[Symbol.dispose]=function(){this.dispose()};H.prototype.H=function(){if(this.g)for(;this.g.length;)this.g.shift()()};var I=function(a,b){this.type=a;this.g=this.target=b;this.defaultPrevented=!1};I.prototype.h=function(){this.defaultPrevented=!0};var Ja=function(){if(!t.addEventListener||!Object.defineProperty)return!1;var a=!1,b=Object.defineProperty({},"passive",{get:function(){a=!0}});try{var c=function(){};t.addEventListener("test",c,b);t.removeEventListener("test",c,b)}catch(d){}return a}();var J=function(a,b){I.call(this,a?a.type:"");this.relatedTarget=this.g=this.target=null;this.button=this.screenY=this.screenX=this.clientY=this.clientX=0;this.key="";this.metaKey=this.shiftKey=this.altKey=this.ctrlKey=!1;this.state=null;this.pointerId=0;this.pointerType="";this.j=null;a&&this.init(a,b)};w(J,I);
J.prototype.init=function(a,b){var c=this.type=a.type,d=a.changedTouches&&a.changedTouches.length?a.changedTouches[0]:null;this.target=a.target||a.srcElement;this.g=b;b=a.relatedTarget;b||(c=="mouseover"?b=a.fromElement:c=="mouseout"&&(b=a.toElement));this.relatedTarget=b;d?(this.clientX=d.clientX!==void 0?d.clientX:d.pageX,this.clientY=d.clientY!==void 0?d.clientY:d.pageY,this.screenX=d.screenX||0,this.screenY=d.screenY||0):(this.clientX=a.clientX!==void 0?a.clientX:a.pageX,this.clientY=a.clientY!==
void 0?a.clientY:a.pageY,this.screenX=a.screenX||0,this.screenY=a.screenY||0);this.button=a.button;this.key=a.key||"";this.ctrlKey=a.ctrlKey;this.altKey=a.altKey;this.shiftKey=a.shiftKey;this.metaKey=a.metaKey;this.pointerId=a.pointerId||0;this.pointerType=a.pointerType;this.state=a.state;this.j=a;a.defaultPrevented&&J.P.h.call(this)};J.prototype.h=function(){J.P.h.call(this);var a=this.j;a.preventDefault?a.preventDefault():a.returnValue=!1};var K="closure_listenable_"+(Math.random()*1E6|0);var Ka=0;var La=function(a,b,c,d,e){this.listener=a;this.proxy=null;this.src=b;this.type=c;this.capture=!!d;this.M=e;this.key=++Ka;this.K=this.L=!1},L=function(a){a.K=!0;a.listener=null;a.proxy=null;a.src=null;a.M=null};var Ma="constructor hasOwnProperty isPrototypeOf propertyIsEnumerable toLocaleString toString valueOf".split(" ");function Na(a,b){for(var c,d,e=1;e<arguments.length;e++){d=arguments[e];for(c in d)a[c]=d[c];for(var f=0;f<Ma.length;f++)c=Ma[f],Object.prototype.hasOwnProperty.call(d,c)&&(a[c]=d[c])}};function M(a){this.src=a;this.g={};this.h=0}M.prototype.add=function(a,b,c,d,e){var f=a.toString();a=this.g[f];a||(a=this.g[f]=[],this.h++);var k=Oa(a,b,d,e);k>-1?(b=a[k],c||(b.L=!1)):(b=new La(b,this.src,f,!!d,e),b.L=c,a.push(b));return b};var Pa=function(a,b){var c=b.type;c in a.g&&sa(a.g[c],b)&&(L(b),a.g[c].length==0&&(delete a.g[c],a.h--))},Oa=function(a,b,c,d){for(var e=0;e<a.length;++e){var f=a[e];if(!f.K&&f.listener==b&&f.capture==!!c&&f.M==d)return e}return-1};var Qa="closure_lm_"+(Math.random()*1E6|0),Ra={},Sa=0,Ua=function(a,b,c,d,e){if(d&&d.once)Ta(a,b,c,d,e);else if(Array.isArray(b))for(var f=0;f<b.length;f++)Ua(a,b[f],c,d,e);else c=Va(c),a&&a[K]?(d=u(d)?!!d.capture:!!d,Wa(a),a.u.add(String(b),c,!1,d,e)):Xa(a,b,c,!1,d,e)},Xa=function(a,b,c,d,e,f){if(!b)throw Error("Invalid event type");var k=u(e)?!!e.capture:!!e,g=Ya(a);g||(a[Qa]=g=new M(a));c=g.add(b,c,d,k,f);if(!c.proxy){d=Za();c.proxy=d;d.src=a;d.listener=c;if(a.addEventListener)Ja||(e=k),e===void 0&&
(e=!1),a.addEventListener(b.toString(),d,e);else if(a.attachEvent)a.attachEvent($a(b.toString()),d);else if(a.addListener&&a.removeListener)A(b==="change","MediaQueryList only has a change event"),a.addListener(d);else throw Error("addEventListener and attachEvent are unavailable.");Sa++}},Za=function(){var a=ab,b=function(c){return a.call(b.src,b.listener,c)};return b},Ta=function(a,b,c,d,e){if(Array.isArray(b))for(var f=0;f<b.length;f++)Ta(a,b[f],c,d,e);else c=Va(c),a&&a[K]?a.u.add(String(b),c,
!0,u(d)?!!d.capture:!!d,e):Xa(a,b,c,!0,d,e)},bb=function(a,b,c,d,e){if(Array.isArray(b))for(var f=0;f<b.length;f++)bb(a,b[f],c,d,e);else(d=u(d)?!!d.capture:!!d,c=Va(c),a&&a[K])?(a=a.u,b=String(b).toString(),b in a.g&&(f=a.g[b],c=Oa(f,c,d,e),c>-1&&(L(f[c]),A(f.length!=null),Array.prototype.splice.call(f,c,1),f.length==0&&(delete a.g[b],a.h--)))):a&&(a=Ya(a))&&(b=a.g[b.toString()],a=-1,b&&(a=Oa(b,c,d,e)),(c=a>-1?b[a]:null)&&cb(c))},cb=function(a){if(typeof a!=="number"&&a&&!a.K){var b=a.src;if(b&&b[K])Pa(b.u,
a);else{var c=a.type,d=a.proxy;b.removeEventListener?b.removeEventListener(c,d,a.capture):b.detachEvent?b.detachEvent($a(c),d):b.addListener&&b.removeListener&&b.removeListener(d);Sa--;(c=Ya(b))?(Pa(c,a),c.h==0&&(c.src=null,b[Qa]=null)):L(a)}}},$a=function(a){return a in Ra?Ra[a]:Ra[a]="on"+a},ab=function(a,b){if(a.K)a=!0;else{b=new J(b,this);var c=a.listener,d=a.M||a.src;a.L&&cb(a);a=c.call(d,b)}return a},Ya=function(a){a=a[Qa];return a instanceof M?a:null},db="__closure_events_fn_"+(Math.random()*
1E9>>>0),Va=function(a){A(a,"Listener can not be null.");if(typeof a==="function")return a;A(a.handleEvent,"An object listener must have handleEvent method.");a[db]||(a[db]=function(b){return a.handleEvent(b)});return a[db]};var N=function(){H.call(this);this.u=new M(this);this.j=this;this.h=null};w(N,H);N.prototype[K]=!0;N.prototype.addEventListener=function(a,b,c,d){Ua(this,a,b,c,d)};N.prototype.removeEventListener=function(a,b,c,d){bb(this,a,b,c,d)};
N.prototype.dispatchEvent=function(a){Wa(this);var b=this.h;if(b){var c=[];for(var d=1;b;b=b.h)c.push(b),A(++d<1E3,"infinite loop")}b=this.j;d=a.type||a;if(typeof a==="string")a=new I(a,b);else if(a instanceof I)a.target=a.target||b;else{var e=a;a=new I(d,b);Na(a,e)}e=!0;var f;if(c)for(f=c.length-1;f>=0;f--){var k=a.g=c[f];e=O(k,d,!0,a)&&e}k=a.g=b;e=O(k,d,!0,a)&&e;e=O(k,d,!1,a)&&e;if(c)for(f=0;f<c.length;f++)k=a.g=c[f],e=O(k,d,!1,a)&&e;return e};
N.prototype.H=function(){N.P.H.call(this);if(this.u){var a=this.u,b=0,c;for(c in a.g){for(var d=a.g[c],e=0;e<d.length;e++)++b,L(d[e]);delete a.g[c];a.h--}}this.h=null};var O=function(a,b,c,d){b=a.u.g[String(b)];if(!b)return!0;b=b.concat();for(var e=!0,f=0;f<b.length;++f){var k=b[f];if(k&&!k.K&&k.capture==c){var g=k.listener,h=k.M||k.src;k.L&&Pa(a.u,k);e=g.call(h,d)!==!1&&e}}return e&&!d.defaultPrevented},Wa=function(a){A(a.u,"Event target is not initialized. Did you call the superclass (goog.events.EventTarget) constructor?")};var eb=RegExp("^(?:([^:/?#.]+):)?(?://(?:([^\\\\/?#]*)@)?([^\\\\/?#]*?)(?::([0-9]+))?(?=[\\\\/?#]|$))?([^?#]+)?(?:\\?([^#]*))?(?:#([\\s\\S]*))?$"),fb=function(a,b){if(a){a=a.split("&");for(var c=0;c<a.length;c++){var d=a[c].indexOf("="),e=null;if(d>=0){var f=a[c].substring(0,d);e=a[c].substring(d+1)}else f=a[c];b(f,e?decodeURIComponent(e.replace(/\+/g," ")):"")}}};var P=function(){N.call(this);this.headers=new Map;this.A=!1;this.i=null;this.J=this.W=this.O="";this.B=this.U=this.N=this.T=!1;this.R=0;this.F=null;this.Z="";this.da=this.aa=!1;this.S=this.V=null};w(P,N);P.prototype.s=E(Fa(),"goog.net.XhrIo").o;var gb=/^https?$/i,hb=["POST","PUT"],ib=[];P.prototype.ba=function(){this.dispose();sa(ib,this)};P.prototype.setTrustToken=function(a){this.V=a};P.prototype.setAttributionReporting=function(a){this.S=a};
P.prototype.send=function(a,b,c,d){if(this.i)throw Error("[goog.net.XhrIo] Object is active with another request="+this.O+"; newUri="+a);b=b?b.toUpperCase():"GET";this.O=a;this.J="";this.W=b;this.T=!1;this.A=!0;this.i=new XMLHttpRequest;this.i.onreadystatechange=Ia(v(this.Y,this));this.da&&"onprogress"in this.i&&(this.i.onprogress=Ia(v(function(k){this.X(k,!0)},this)),this.i.upload&&(this.i.upload.onprogress=Ia(v(this.X,this))));try{F(this.s,Q(this,"Opening Xhr")),this.U=!0,this.i.open(b,String(a),
!0),this.U=!1}catch(k){F(this.s,Q(this,"Error opening Xhr: "+k.message));jb(this,k);return}a=c||"";c=new Map(this.headers);if(d)if(Object.getPrototypeOf(d)===Object.prototype)for(var e in d)c.set(e,d[e]);else if(typeof d.keys==="function"&&typeof d.get==="function"){e=q(d.keys());for(var f=e.next();!f.done;f=e.next())f=f.value,c.set(f,d.get(f))}else throw Error("Unknown input type for opt_headers: "+String(d));d=Array.from(c.keys()).find(function(k){return"content-type"==k.toLowerCase()});e=t.FormData&&
a instanceof t.FormData;!(ra(hb,b)>=0)||d||e||c.set("Content-Type","application/x-www-form-urlencoded;charset=utf-8");b=q(c);for(d=b.next();!d.done;d=b.next())c=q(d.value),d=c.next().value,c=c.next().value,this.i.setRequestHeader(d,c);this.Z&&(this.i.responseType=this.Z);"withCredentials"in this.i&&this.i.withCredentials!==this.aa&&(this.i.withCredentials=this.aa);if("setTrustToken"in this.i&&this.V)try{this.i.setTrustToken(this.V)}catch(k){F(this.s,Q(this,"Error SetTrustToken: "+k.message))}if("setAttributionReporting"in
this.i&&this.S)try{this.i.setAttributionReporting(this.S)}catch(k){F(this.s,Q(this,"Error SetAttributionReporting: "+k.message))}try{this.F&&(clearTimeout(this.F),this.F=null),this.R>0&&(F(this.s,Q(this,"Will abort after "+this.R+"ms if incomplete")),this.F=setTimeout(this.ea.bind(this),this.R)),F(this.s,Q(this,"Sending request")),this.N=!0,this.i.send(a),this.N=!1}catch(k){F(this.s,Q(this,"Send error: "+k.message)),jb(this,k)}};
P.prototype.ea=function(){typeof fa!="undefined"&&this.i&&(this.J="Timed out after "+this.R+"ms, aborting",F(this.s,Q(this,this.J)),this.dispatchEvent("timeout"),this.abort(8))};var jb=function(a,b){a.A=!1;a.i&&(a.B=!0,a.i.abort(),a.B=!1);a.J=b;kb(a);R(a)},kb=function(a){a.T||(a.T=!0,a.dispatchEvent("complete"),a.dispatchEvent("error"))};
P.prototype.abort=function(){this.i&&this.A&&(F(this.s,Q(this,"Aborting")),this.A=!1,this.B=!0,this.i.abort(),this.B=!1,this.dispatchEvent("complete"),this.dispatchEvent("abort"),R(this))};P.prototype.H=function(){this.i&&(this.A&&(this.A=!1,this.B=!0,this.i.abort(),this.B=!1),R(this,!0));P.P.H.call(this)};P.prototype.Y=function(){this.I||(this.U||this.N||this.B?lb(this):this.ca())};P.prototype.ca=function(){lb(this)};
var lb=function(a){if(a.A&&typeof fa!="undefined")if(a.N&&S(a)==4)setTimeout(a.Y.bind(a),0);else if(a.dispatchEvent("readystatechange"),S(a)==4){F(a.s,Q(a,"Request complete"));a.A=!1;try{if(mb(a))a.dispatchEvent("complete"),a.dispatchEvent("success");else{try{var b=S(a)>2?a.i.statusText:""}catch(c){F(a.s,"Can not get status: "+c.message),b=""}a.J=b+" ["+nb(a)+"]";kb(a)}}finally{R(a)}}};
P.prototype.X=function(a,b){A(a.type==="progress","goog.net.EventType.PROGRESS is of the same type as raw XHR progress.");this.dispatchEvent(ob(a,"progress"));this.dispatchEvent(ob(a,b?"downloadprogress":"uploadprogress"))};
var ob=function(a,b){return{type:b,lengthComputable:a.lengthComputable,loaded:a.loaded,total:a.total}},R=function(a,b){if(a.i){a.F&&(clearTimeout(a.F),a.F=null);var c=a.i;a.i=null;b||a.dispatchEvent("ready");try{c.onreadystatechange=null}catch(d){(a=a.s)&&Ga(a,ua,"Problem encountered resetting onreadystatechange: "+d.message)}}};P.prototype.isActive=function(){return!!this.i};
var mb=function(a){var b=nb(a);a:switch(b){case 200:case 201:case 202:case 204:case 206:case 304:case 1223:var c=!0;break a;default:c=!1}if(!c){if(b=b===0)a=String(a.O).match(eb)[1]||null,!a&&t.self&&t.self.location&&(a=t.self.location.protocol.slice(0,-1)),b=!gb.test(a?a.toLowerCase():"");c=b}return c},S=function(a){return a.i?a.i.readyState:0},nb=function(a){try{return S(a)>2?a.i.status:-1}catch(b){return-1}};
P.prototype.getResponseHeader=function(a){if(this.i&&S(this)==4)return a=this.i.getResponseHeader(a),a===null?void 0:a};P.prototype.getAllResponseHeaders=function(){return this.i&&S(this)>=2?this.i.getAllResponseHeaders()||"":""};var Q=function(a,b){return b+" ["+a.W+" "+a.O+" "+nb(a)+"]"};var T=function(a){this.g=this.D=this.l="";this.G=null;this.C=this.h="";this.o=!1;var b;a instanceof T?(this.o=a.o,pb(this,a.l),this.D=a.D,this.g=a.g,qb(this,a.G),U(this,a.h),rb(this,sb(a.j)),this.C=a.C):a&&(b=String(a).match(eb))?(this.o=!1,pb(this,b[1]||"",!0),this.D=V(b[2]||""),this.g=V(b[3]||"",!0),qb(this,b[4]),U(this,b[5]||"",!0),rb(this,b[6]||"",!0),this.C=V(b[7]||"")):(this.o=!1,this.j=new W(null,this.o))};
T.prototype.toString=function(){var a=[],b=this.l;b&&a.push(X(b,tb,!0),":");var c=this.g;if(c||b=="file")a.push("//"),(b=this.D)&&a.push(X(b,tb,!0),"@"),a.push(encodeURIComponent(String(c)).replace(/%25([0-9a-fA-F]{2})/g,"%$1")),c=this.G,c!=null&&a.push(":",String(c));if(c=this.h)this.g&&c.charAt(0)!="/"&&a.push("/"),a.push(X(c,c.charAt(0)=="/"?ub:vb,!0));(c=this.j.toString())&&a.push("?",c);(c=this.C)&&a.push("#",X(c,wb));return a.join("")};
T.prototype.resolve=function(a){var b=new T(this),c=!!a.l;c?pb(b,a.l):c=!!a.D;c?b.D=a.D:c=!!a.g;c?b.g=a.g:c=a.G!=null;var d=a.h;if(c)qb(b,a.G);else if(c=!!a.h){if(d.charAt(0)!="/")if(this.g&&!this.h)d="/"+d;else{var e=b.h.lastIndexOf("/");e!=-1&&(d=b.h.slice(0,e+1)+d)}e=d;if(e==".."||e==".")d="";else if(e.indexOf("./")!=-1||e.indexOf("/.")!=-1){d=e.lastIndexOf("/",0)==0;e=e.split("/");for(var f=[],k=0;k<e.length;){var g=e[k++];g=="."?d&&k==e.length&&f.push(""):g==".."?((f.length>1||f.length==1&&f[0]!=
"")&&f.pop(),d&&k==e.length&&f.push("")):(f.push(g),d=!0)}d=f.join("/")}else d=e}c?U(b,d):c=a.j.toString()!=="";c?rb(b,sb(a.j)):c=!!a.C;c&&(b.C=a.C);return b};
var pb=function(a,b,c){a.l=c?V(b,!0):b;a.l&&(a.l=a.l.replace(/:$/,""))},qb=function(a,b){if(b){b=Number(b);if(isNaN(b)||b<0)throw Error("Bad port number "+b);a.G=b}else a.G=null},U=function(a,b,c){a.h=c?V(b,!0):b;return a},rb=function(a,b,c){b instanceof W?(a.j=b,xb(a.j,a.o)):(c||(b=X(b,yb)),a.j=new W(b,a.o));return a},V=function(a,b){return a?b?decodeURI(a.replace(/%25/g,"%2525")):decodeURIComponent(a):""},X=function(a,b,c){return typeof a==="string"?(a=encodeURI(a).replace(b,zb),c&&(a=a.replace(/%25([0-9a-fA-F]{2})/g,
"%$1")),a):null},zb=function(a){a=a.charCodeAt(0);return"%"+(a>>4&15).toString(16)+(a&15).toString(16)},tb=/[#\/\?@]/g,vb=/[#\?:]/g,ub=/[#\?]/g,yb=/[#\?@]/g,wb=/#/g,W=function(a,b){this.h=this.g=null;this.j=a||null;this.l=!!b},Y=function(a){a.g||(a.g=new Map,a.h=0,a.j&&fb(a.j,function(b,c){a.add(decodeURIComponent(b.replace(/\+/g," ")),c)}))};W.prototype.add=function(a,b){Y(this);this.j=null;a=Z(this,a);var c=this.g.get(a);c||this.g.set(a,c=[]);c.push(b);this.h=C(this.h)+1;return this};
var Ab=function(a,b){Y(a);b=Z(a,b);a.g.has(b)&&(a.j=null,a.h=C(a.h)-a.g.get(b).length,a.g.delete(b))},Bb=function(a,b){Y(a);b=Z(a,b);return a.g.has(b)};W.prototype.forEach=function(a,b){Y(this);this.g.forEach(function(c,d){c.forEach(function(e){a.call(b,e,d,this)},this)},this)};W.prototype.o=function(a){Y(this);var b=[];if(typeof a==="string")Bb(this,a)&&(b=b.concat(this.g.get(Z(this,a))));else{a=Array.from(this.g.values());for(var c=0;c<a.length;c++)b=b.concat(a[c])}return b};
W.prototype.set=function(a,b){Y(this);this.j=null;a=Z(this,a);Bb(this,a)&&(this.h=C(this.h)-this.g.get(a).length);this.g.set(a,[b]);this.h=C(this.h)+1;return this};W.prototype.get=function(a,b){if(!a)return b;a=this.o(a);return a.length>0?String(a[0]):b};
W.prototype.toString=function(){if(this.j)return this.j;if(!this.g)return"";for(var a=[],b=Array.from(this.g.keys()),c=0;c<b.length;c++){var d=b[c],e=encodeURIComponent(String(d));d=this.o(d);for(var f=0;f<d.length;f++){var k=e;d[f]!==""&&(k+="="+encodeURIComponent(String(d[f])));a.push(k)}}return this.j=a.join("&")};
var sb=function(a){var b=new W;b.j=a.j;a.g&&(b.g=new Map(a.g),b.h=a.h);return b},Z=function(a,b){b=String(b);a.l&&(b=b.toLowerCase());return b},xb=function(a,b){b&&!a.l&&(Y(a),a.j=null,a.g.forEach(function(c,d){var e=d.toLowerCase();if(d!=e&&(Ab(this,d),Ab(this,e),c.length>0)){this.j=null;d=this.g;var f=d.set;e=Z(this,e);var k=c.length;if(k>0){for(var g=Array(k),h=0;h<k;h++)g[h]=c[h];k=g}else k=[];f.call(d,e,k);this.h=C(this.h)+c.length}},a));a.l=b};var Db=function(){this.h=void 0;this.g=null;Cb(this,0);window.addEventListener("load",this.o.bind(this))};
Db.prototype.l=function(a){if(this.g){a=a.target;var b;if(b=mb(a)){try{var c=a.i?a.i.responseText:""}catch(d){F(a.s,"Can not get responseText: "+d.message),c=""}b=c==="OK"}if(b){this.j();c=window.location;a=U(new T(window.location),"/ServiceLogin").toString();if(a instanceof x)if(a instanceof x)a=a.g;else throw Error("Unexpected type when unwrapping SafeUrl, got '"+a+"' of type '"+typeof a+"'");else(b=!la.test(a))&&na(a),a=b?void 0:a;a!==void 0&&(c.href=a)}else Cb(this,5E3)}};
var Cb=function(a,b){a.g=setTimeout(function(){if(a.g){var c=Ha.get("APISID");if(c===a.h)Cb(a,5E3);else{a.h=c;c=new T("/PassiveLoginProber");var d=(new T(window.location)).j;c=rb(c,d).toString();d=a.l.bind(a);var e=new P;ib.push(e);d&&(Wa(e),e.u.add("complete",d,!1,void 0,void 0));e.u.add("ready",e.ba,!0,void 0,void 0);e.send(c,void 0,void 0,void 0)}}},b)};Db.prototype.o=function(){document.addEventListener("submit",this.j.bind(this))};
Db.prototype.j=function(){this.g&&(clearTimeout(this.g),this.g=null)};new Db;}).call(this);
</script><c-data id="i3"></c-data></c-wiz></div></section></div><span jsslot><div class="D4rY0b"><p class="vOZun">Not your computer? Use a private browsing window to sign in. <a href="https://support.google.com/accounts?p=signin_privatebrowsing&amp;hl=en-US" jsname="JFyozc" target="_blank">Learn more about using Guest mode</a></p></div></span><div class="i2knIc" jsname="DH6Rkf"><div class="wg0fFb" jsname="DhK0U"><div class="RhTxBf" jsname="k77Iif"><button name="action" class="JnOM6e TrZEUc rDisVe" value="1" jsname="Njthtb" id="identifierNext">Next</button></div><div class="tmMcIf" jsname="QkNstf"><a href="/lifecycle/flows/signup?continue=https://drive.usercontent.google.com/download?id%3D15vEesL8xTMFSo-uLA5dsx3puVaKcGEyw%26export%3Ddownload&amp;dsh=S707491678:1743896408202977&amp;flowEntry=SignUp&amp;flowName=GlifWebSignIn&amp;followup=https://drive.usercontent.google.com/download?id%3D15vEesL8xTMFSo-uLA5dsx3puVaKcGEyw%26export%3Ddownload&amp;ifkv=AXH0vVv0CbiU_Wk9REDVCw4rixpQn-GDo7--KsMDAK3yiLZzH0XMmVwFpBv9kkMWTOzwD-UHys9d&amp;service=wise" class="JnOM6e TrZEUc kTeh9 KXbQ4b">Create account</a></div></div></div><input type="hidden" name="at" value="AAQ76x6_JXCw8bmV_VwGxSai1Odh:1743896408304"></form></div></div><script aria-hidden="true" nonce="c6XQoK_6ljSIPUPPhVJTog">window.wiz_progress&&window.wiz_progress();window.wiz_tick&&window.wiz_tick('chA7fe');</script></body></html></div><c-wiz jsrenderer="ZdRp7e" jsshadow jsdata="deferred-i1" data-node-index="0;0" jsmodel="hc6Ubd" c-wiz><footer class="HUYFt" data-auto-init="Footer"><div class="hXs2T"><form autocomplete="off"><select name="hl" class="N158t" data-language-selector-select jsname="rfCUpd"><option value="af">Afrikaans</option><option value="az">azərbaycan</option><option value="bs">bosanski</option><option value="ca">català</option><option value="cs">Čeština</option><option value="cy">Cymraeg</option><option value="da">Dansk</option><option value="de">Deutsch</option><option value="et">eesti</option><option value="en-GB">English (United Kingdom)</option><option value="en-US" selected>English (United States)</option><option value="es-ES">Español (España)</option><option value="es-419">Español (Latinoamérica)</option><option value="eu">euskara</option><option value="fil">Filipino</option><option value="fr-CA">Français (Canada)</option><option value="fr-FR">Français (France)</option><option value="ga">Gaeilge</option><option value="gl">galego</option><option value="hr">Hrvatski</option><option value="id">Indonesia</option><option value="zu">isiZulu</option><option value="is">íslenska</option><option value="it">Italiano</option><option value="sw">Kiswahili</option><option value="lv">latviešu</option><option value="lt">lietuvių</option><option value="hu">magyar</option><option value="ms">Melayu</option><option value="nl">Nederlands</option><option value="no">norsk</option><option value="uz">o‘zbek</option><option value="pl">polski</option><option value="pt-BR">Português (Brasil)</option><option value="pt-PT">Português (Portugal)</option><option value="ro">română</option><option value="sq">shqip</option><option value="sk">Slovenčina</option><option value="sl">slovenščina</option><option value="sr-Latn">srpski (latinica)</option><option value="fi">Suomi</option><option value="sv">Svenska</option><option value="vi">Tiếng Việt</option><option value="tr">Türkçe</option><option value="el">Ελληνικά</option><option value="be">беларуская</option><option value="bg">български</option><option value="ky">кыргызча</option><option value="kk">қазақ тілі</option><option value="mk">македонски</option><option value="mn">монгол</option><option value="ru">Русский</option><option value="sr-Cyrl">српски (ћирилица)</option><option value="uk">Українська</option><option value="ka">ქართული</option><option value="hy">հայերեն</option><option value="iw">‫עברית‬‎</option><option value="ur">‫اردو‬‎</option><option value="ar">‫العربية‬‎</option><option value="fa">‫فارسی‬‎</option><option value="am">አማርኛ</option><option value="ne">नेपाली</option><option value="mr">मराठी</option><option value="hi">हिन्दी</option><option value="as">অসমীয়া</option><option value="bn">বাংলা</option><option value="pa">ਪੰਜਾਬੀ</option><option value="gu">ગુજરાતી</option><option value="or">ଓଡ଼ିଆ</option><option value="ta">தமிழ்</option><option value="te">తెలుగు</option><option value="kn">ಕನ್ನಡ</option><option value="ml">മലയാളം</option><option value="si">සිංහල</option><option value="th">ไทย</option><option value="lo">ລາວ</option><option value="my">မြန်မာ</option><option value="km">ខ្មែរ</option><option value="ko">한국어</option><option value="zh-HK">中文（香港）</option><option value="ja">日本語</option><option value="zh-CN">简体中文</option><option value="zh-TW">繁體中文</option></select></form></div><ul class="M2nKge"><li class="vomtoe"><a class="pUP0Nd TrZEUc" href="https://support.google.com/accounts?hl=en-US&amp;p=account_iph" target="_blank"><span class="UskCyf">Help</span></a></li><li class="vomtoe"><a class="pUP0Nd TrZEUc" href="https://accounts.google.com/TOS?loc=US&amp;hl=en-US&amp;privacy=true" target="_blank"><span class="UskCyf">Privacy</span></a></li><li class="vomtoe"><a class="pUP0Nd TrZEUc" href="https://accounts.google.com/TOS?loc=US&amp;hl=en-US" target="_blank"><span class="UskCyf">Terms</span></a></li></ul></footer><c-data id="i1" jsdata=" OsjLy;_;2"></c-data></c-wiz><script aria-hidden="true" nonce="c6XQoK_6ljSIPUPPhVJTog">window.wiz_progress&&window.wiz_progress();window.wiz_tick&&window.wiz_tick('ZdRp7e');</script><script nonce="c6XQoK_6ljSIPUPPhVJTog">(function(){'use strict';var a=function(b){var c=0;return function(){return c<b.length?{done:!1,value:b[c++]}:{done:!0}}},h=typeof Object.defineProperties=="function"?Object.defineProperty:function(b,c,d){if(b==Array.prototype||b==Object.prototype)return b;b[c]=d.value;return b},aa=function(b){b=["object"==typeof globalThis&&globalThis,b,"object"==typeof window&&window,"object"==typeof self&&self,"object"==typeof global&&global];for(var c=0;c<b.length;++c){var d=b[c];if(d&&d.Math==Math)return d}throw Error("Cannot find global object");
},l=aa(this),m=function(b,c){if(c)a:{var d=l;b=b.split(".");for(var e=0;e<b.length-1;e++){var f=b[e];if(!(f in d))break a;d=d[f]}b=b[b.length-1];e=d[b];c=c(e);c!=e&&c!=null&&h(d,b,{configurable:!0,writable:!0,value:c})}};
m("Symbol",function(b){if(b)return b;var c=function(g,k){this.i=g;h(this,"description",{configurable:!0,writable:!0,value:k})};c.prototype.toString=function(){return this.i};var d="jscomp_symbol_"+(Math.random()*1E9>>>0)+"_",e=0,f=function(g){if(this instanceof f)throw new TypeError("Symbol is not a constructor");return new c(d+(g||"")+"_"+e++,g)};return f});
m("Symbol.iterator",function(b){if(b)return b;b=Symbol("Symbol.iterator");for(var c="Array Int8Array Uint8Array Uint8ClampedArray Int16Array Uint16Array Int32Array Uint32Array Float32Array Float64Array".split(" "),d=0;d<c.length;d++){var e=l[c[d]];typeof e==="function"&&typeof e.prototype[b]!="function"&&h(e.prototype,b,{configurable:!0,writable:!0,value:function(){return ba(a(this))}})}return b});
var ba=function(b){b={next:b};b[Symbol.iterator]=function(){return this};return b},ca=typeof Object.create=="function"?Object.create:function(b){var c=function(){};c.prototype=b;return new c},p;if(typeof Object.setPrototypeOf=="function")p=Object.setPrototypeOf;else{var q;a:{var da={a:!0},r={};try{r.__proto__=da;q=r.a;break a}catch(b){}q=!1}p=q?function(b,c){b.__proto__=c;if(b.__proto__!==c)throw new TypeError(b+" is not extensible");return b}:null}
var u=p,v=function(b,c){b.prototype=ca(c.prototype);b.prototype.constructor=b;if(u)u(b,c);else for(var d in c)if(d!="prototype")if(Object.defineProperties){var e=Object.getOwnPropertyDescriptor(c,d);e&&Object.defineProperty(b,d,e)}else b[d]=c[d];b.o=c.prototype},w=function(b){var c=typeof Symbol!="undefined"&&Symbol.iterator&&b[Symbol.iterator];if(c)return c.call(b);if(typeof b.length=="number")return{next:a(b)};throw Error(String(b)+" is not an iterable or ArrayLike");},ea=function(b){if(!(b instanceof
Array)){b=w(b);for(var c,d=[];!(c=b.next()).done;)d.push(c.value);b=d}return b};m("globalThis",function(b){return b||l});var fa=function(b,c){b instanceof String&&(b+="");var d=0,e=!1,f={next:function(){if(!e&&d<b.length){var g=d++;return{value:c(g,b[g]),done:!1}}e=!0;return{done:!0,value:void 0}}};f[Symbol.iterator]=function(){return f};return f};m("Array.prototype.keys",function(b){return b?b:function(){return fa(this,function(c){return c})}});/*

 Copyright The Closure Library Authors.
 SPDX-License-Identifier: Apache-2.0
*/
var x=function(b,c){function d(){}d.prototype=c.prototype;b.o=c.prototype;b.prototype=new d;b.prototype.constructor=b;b.s=function(e,f,g){for(var k=Array(arguments.length-2),n=2;n<arguments.length;n++)k[n-2]=arguments[n];return c.prototype[f].apply(e,k)}};var y=function(b){this.i=b;this.l()};function z(b,c){if(Error.captureStackTrace)Error.captureStackTrace(this,z);else{var d=Error().stack;d&&(this.stack=d)}b&&(this.message=String(b));c!==void 0&&(this.cause=c)}x(z,Error);z.prototype.name="CustomError";function A(b,c){b=b.split("%s");for(var d="",e=b.length-1,f=0;f<e;f++)d+=b[f]+(f<c.length?c[f]:"%s");z.call(this,d+b[e])}x(A,z);A.prototype.name="AssertionError";var B=function(b,c,d){if(!b){var e="Assertion failed";if(c){e+=": "+c;var f=Array.prototype.slice.call(arguments,2)}throw new A(""+e,f||[]);}return b};var C=function(){y.apply(this,arguments);this.j=!1};v(C,y);C.prototype.l=function(){var b=this;this.j=this.i.dataset.isRemoveMode==="true";var c;(c=this.i.querySelector("[data-rab]"))==null||c.addEventListener("click",function(e){e.preventDefault();D(b,!0)});var d;(d=this.i.querySelector("[data-radb]"))==null||d.addEventListener("click",function(e){e.preventDefault();D(b,!1)})};
var D=function(b,c){b.j!==c&&(b.j=c,b.i.dataset.isRemoveMode=c.toString(),b.i.querySelectorAll("[data-ci]").forEach(function(d){d.getElementsByTagName("BUTTON".toString()).item(0).name=b.j?"chooser[remove]":"chooser[select]"}))};var E=function(){y.apply(this,arguments)};v(E,y);E.prototype.l=function(){var b=this.i.querySelector("FORM".toString());b&&this.i.addEventListener("submit",function(c){b.getAttribute("data-is-submitted")==="true"?c.preventDefault():b.setAttribute("data-is-submitted","true")})};/*

 Copyright Google LLC
 SPDX-License-Identifier: Apache-2.0
*/
var F={};function G(){if(F!==F)throw Error("Bad secret");};var H=globalThis.trustedTypes,I;function ha(){var b=null;if(!H)return b;try{var c=function(d){return d};b=H.createPolicy("goog#html",{createHTML:c,createScript:c,createScriptURL:c})}catch(d){throw d;}return b};var J=function(b){G();this.i=b};J.prototype.toString=function(){return this.i};new J("about:blank");new J("about:invalid#zClosurez");var ia=/^\s*(?!javascript:)(?:[\w+.-]+:|[^:/?#]*(?:[/?#]|$))/i,K=[],L=function(){};ja(function(b){console.warn("A URL with content '"+b+"' was sanitized away.")});function ja(b){K.indexOf(b)===-1&&K.push(b);L=function(c){K.forEach(function(d){d(c)})}};var M=function(b){G();this.i=b};M.prototype.toString=function(){return this.i+""};var N=function(){y.apply(this,arguments)};v(N,y);N.prototype.l=function(){var b=this.i.querySelector("[data-language-selector-select]");b&&ka(b)};
function ka(b){b.addEventListener("change",function(c){c=c.target;if(c.value){var d=new URL(document.location.toString());d.searchParams.set("hl",c.value);c=window.location;d=d.toString();if(d instanceof J)if(d instanceof J)d=d.i;else throw Error("Unexpected type when unwrapping SafeUrl, got '"+d+"' of type '"+typeof d+"'");else{var e=!ia.test(d);e&&L(d);d=e?void 0:d}d!==void 0&&(c.href=d)}})};var O=Object.create(null);function P(b,c){O[b]||(O[b]=c)};var Q=function(){y.apply(this,arguments)};v(Q,y);Q.prototype.l=function(){var b=this.i.querySelector("#playCaptchaButton"),c=this.i.querySelector("#captchaAudio"),d=this.i.querySelector("input[name=ca]");b&&c&&d&&b.addEventListener("click",function(e){e.preventDefault();c.readyState===HTMLMediaElement.HAVE_NOTHING?c.load():c.paused&&c.play();d.value="";d.focus()})};var R=function(){y.apply(this,arguments)};v(R,y);R.prototype.l=function(){this.i.dataset.hasDomainSuffix!==void 0&&(S(this.i),la(this.i))};function la(b){b.addEventListener("keyup",function(){S(b)})}function S(b){b.getElementsByTagName("INPUT".toString()).item(0).value.indexOf("@")>0?b.dataset.hasAtSign="":delete b.dataset.hasAtSign};var T=function(){y.apply(this,arguments);this.j=0};v(T,y);T.prototype.l=function(){var b=this,c=B(this.i.querySelector("[jsname='Mi0fJc']")).id,d=B(this.i.dataset.siteKey);window.grecaptcha.ready(function(){ma(b,d,c)})};var ma=function(b,c,d){b.j=window.grecaptcha.render(d,{sitekey:c,callback:function(e){B(b.i.querySelector("[jsname='BhKThb']")).setAttribute("value",e)},"expired-callback":function(){window.grecaptcha.reset(b.j)}})};var U=function(){y.apply(this,arguments)};v(U,y);U.prototype.l=function(){var b=this.i;b.dataset.hasDomainSuffix!==void 0&&(na(b),oa(b))};function oa(b){b.addEventListener("keyup",function(){na(b)})}function na(b){b.getElementsByTagName("INPUT".toString()).item(0).value.indexOf("@")>0?b.dataset.hasAtSign="":delete b.dataset.hasAtSign};var V={COUNTRY:{"001":"world","002":"Africa","003":"North America","005":"South America","009":"Oceania","011":"Western Africa","013":"Central America","014":"Eastern Africa","015":"Northern Africa","017":"Middle Africa","018":"Southern Africa","019":"Americas","021":"Northern America","029":"Caribbean","030":"Eastern Asia","034":"Southern Asia","035":"Southeast Asia","039":"Southern Europe","053":"Australasia","054":"Melanesia","057":"Micronesian Region","061":"Polynesia",142:"Asia",143:"Central Asia",
145:"Western Asia",150:"Europe",151:"Eastern Europe",154:"Northern Europe",155:"Western Europe",202:"Sub-Saharan Africa",419:"Latin America",AC:"Ascension Island",AD:"Andorra",AE:"United Arab Emirates",AF:"Afghanistan",AG:"Antigua & Barbuda",AI:"Anguilla",AL:"Albania",AM:"Armenia",AO:"Angola",AQ:"Antarctica",AR:"Argentina",AS:"American Samoa",AT:"Austria",AU:"Australia",AW:"Aruba",AX:"\u00c5land Islands",AZ:"Azerbaijan",BA:"Bosnia & Herzegovina",BB:"Barbados",BD:"Bangladesh",BE:"Belgium",BF:"Burkina Faso",
BG:"Bulgaria",BH:"Bahrain",BI:"Burundi",BJ:"Benin",BL:"St. Barth\u00e9lemy",BM:"Bermuda",BN:"Brunei",BO:"Bolivia",BQ:"Caribbean Netherlands",BR:"Brazil",BS:"Bahamas",BT:"Bhutan",BV:"Bouvet Island",BW:"Botswana",BY:"Belarus",BZ:"Belize",CA:"Canada",CC:"Cocos (Keeling) Islands",CD:"Congo - Kinshasa",CF:"Central African Republic",CG:"Congo - Brazzaville",CH:"Switzerland",CI:"C\u00f4te d\u2019Ivoire",CK:"Cook Islands",CL:"Chile",CM:"Cameroon",CN:"China",CO:"Colombia",CP:"Clipperton Island",CQ:"Sark",
CR:"Costa Rica",CU:"Cuba",CV:"Cape Verde",CW:"Cura\u00e7ao",CX:"Christmas Island",CY:"Cyprus",CZ:"Czechia",DE:"Germany",DG:"Diego Garcia",DJ:"Djibouti",DK:"Denmark",DM:"Dominica",DO:"Dominican Republic",DZ:"Algeria",EA:"Ceuta & Melilla",EC:"Ecuador",EE:"Estonia",EG:"Egypt",EH:"Western Sahara",ER:"Eritrea",ES:"Spain",ET:"Ethiopia",EU:"European Union",EZ:"Eurozone",FI:"Finland",FJ:"Fiji",FK:"Falkland Islands (Islas Malvinas)",FM:"Micronesia",FO:"Faroe Islands",FR:"France",GA:"Gabon",GB:"United Kingdom",
GD:"Grenada",GE:"Georgia",GF:"French Guiana",GG:"Guernsey",GH:"Ghana",GI:"Gibraltar",GL:"Greenland",GM:"Gambia",GN:"Guinea",GP:"Guadeloupe",GQ:"Equatorial Guinea",GR:"Greece",GS:"South Georgia & South Sandwich Islands",GT:"Guatemala",GU:"Guam",GW:"Guinea-Bissau",GY:"Guyana",HK:"Hong Kong",HM:"Heard & McDonald Islands",HN:"Honduras",HR:"Croatia",HT:"Haiti",HU:"Hungary",IC:"Canary Islands",ID:"Indonesia",IE:"Ireland",IL:"Israel",IM:"Isle of Man",IN:"India",IO:"British Indian Ocean Territory",IQ:"Iraq",
IR:"Iran",IS:"Iceland",IT:"Italy",JE:"Jersey",JM:"Jamaica",JO:"Jordan",JP:"Japan",KE:"Kenya",KG:"Kyrgyzstan",KH:"Cambodia",KI:"Kiribati",KM:"Comoros",KN:"St. Kitts & Nevis",KP:"North Korea",KR:"South Korea",KW:"Kuwait",KY:"Cayman Islands",KZ:"Kazakhstan",LA:"Laos",LB:"Lebanon",LC:"St. Lucia",LI:"Liechtenstein",LK:"Sri Lanka",LR:"Liberia",LS:"Lesotho",LT:"Lithuania",LU:"Luxembourg",LV:"Latvia",LY:"Libya",MA:"Morocco",MC:"Monaco",MD:"Moldova",ME:"Montenegro",MF:"St. Martin",MG:"Madagascar",MH:"Marshall Islands",
MK:"North Macedonia",ML:"Mali",MM:"Myanmar (Burma)",MN:"Mongolia",MO:"Macao",MP:"Northern Mariana Islands",MQ:"Martinique",MR:"Mauritania",MS:"Montserrat",MT:"Malta",MU:"Mauritius",MV:"Maldives",MW:"Malawi",MX:"Mexico",MY:"Malaysia",MZ:"Mozambique",NA:"Namibia",NC:"New Caledonia",NE:"Niger",NF:"Norfolk Island",NG:"Nigeria",NI:"Nicaragua",NL:"Netherlands",NO:"Norway",NP:"Nepal",NR:"Nauru",NU:"Niue",NZ:"New Zealand",OM:"Oman",PA:"Panama",PE:"Peru",PF:"French Polynesia",PG:"Papua New Guinea",PH:"Philippines",
PK:"Pakistan",PL:"Poland",PM:"St. Pierre & Miquelon",PN:"Pitcairn Islands",PR:"Puerto Rico",PS:"Palestine",PT:"Portugal",PW:"Palau",PY:"Paraguay",QA:"Qatar",QO:"Outlying Oceania",RE:"R\u00e9union",RO:"Romania",RS:"Serbia",RU:"Russia",RW:"Rwanda",SA:"Saudi Arabia",SB:"Solomon Islands",SC:"Seychelles",SD:"Sudan",SE:"Sweden",SG:"Singapore",SH:"St. Helena",SI:"Slovenia",SJ:"Svalbard & Jan Mayen",SK:"Slovakia",SL:"Sierra Leone",SM:"San Marino",SN:"Senegal",SO:"Somalia",SR:"Suriname",SS:"South Sudan",ST:"S\u00e3o Tom\u00e9 & Pr\u00edncipe",
SV:"El Salvador",SX:"Sint Maarten",SY:"Syria",SZ:"Eswatini",TA:"Tristan da Cunha",TC:"Turks & Caicos Islands",TD:"Chad",TF:"French Southern Territories",TG:"Togo",TH:"Thailand",TJ:"Tajikistan",TK:"Tokelau",TL:"Timor-Leste",TM:"Turkmenistan",TN:"Tunisia",TO:"Tonga",TR:"T\u00fcrkiye",TT:"Trinidad & Tobago",TV:"Tuvalu",TW:"Taiwan",TZ:"Tanzania",UA:"Ukraine",UG:"Uganda",UM:"U.S. Outlying Islands",UN:"United Nations",US:"United States",UY:"Uruguay",UZ:"Uzbekistan",VA:"Vatican City",VC:"St. Vincent & Grenadines",
VE:"Venezuela",VG:"British Virgin Islands",VI:"U.S. Virgin Islands",VN:"Vietnam",VU:"Vanuatu",WF:"Wallis & Futuna",WS:"Samoa",XK:"Kosovo",YE:"Yemen",YT:"Mayotte",ZA:"South Africa",ZM:"Zambia",ZW:"Zimbabwe",ZZ:"Unknown Region"}};var pa={ac:{name:V.COUNTRY.AC,g:"247",index:5},ad:{name:V.COUNTRY.AD,g:"376",index:45},ae:{name:V.COUNTRY.AE,g:"971",index:180},af:{name:V.COUNTRY.AF,g:"93",index:187},ag:{name:V.COUNTRY.AG,g:"1",index:67,h:!0},ai:{name:V.COUNTRY.AI,g:"1",index:158,h:!0},al:{name:V.COUNTRY.AL,g:"355",index:77},am:{name:V.COUNTRY.AM,g:"374",index:12},ao:{name:V.COUNTRY.AO,g:"244",index:155},ar:{name:V.COUNTRY.AR,g:"54",index:193},as:{name:V.COUNTRY.AS,g:"1",index:121,h:!0},at:{name:V.COUNTRY.AT,g:"43",index:102},au:{name:V.COUNTRY.AU,
g:"61",index:134},aw:{name:V.COUNTRY.AW,g:"297",index:60},ax:{name:V.COUNTRY.AX,g:"358",index:235,h:!0},az:{name:V.COUNTRY.AZ,g:"994",index:94},ba:{name:V.COUNTRY.BA,g:"387",index:123},bb:{name:V.COUNTRY.BB,g:"1",index:122,h:!0},bd:{name:V.COUNTRY.BD,g:"880",index:139},be:{name:V.COUNTRY.BE,g:"32",index:0},bf:{name:V.COUNTRY.BF,g:"226",index:56},bg:{name:V.COUNTRY.BG,g:"359",index:208},bh:{name:V.COUNTRY.BH,g:"973",index:115},bi:{name:V.COUNTRY.BI,g:"257",index:150},bj:{name:V.COUNTRY.BJ,g:"229",
index:99},bl:{name:V.COUNTRY.BL,g:"590",index:19,h:!0},bm:{name:V.COUNTRY.BM,g:"1",index:152,h:!0},bn:{name:V.COUNTRY.BN,g:"673",index:131},bo:{name:V.COUNTRY.BO,g:"591",index:128},bq:{name:V.COUNTRY.BQ,g:"599",index:220,h:!0},br:{name:V.COUNTRY.BR,g:"55",index:59},bs:{name:V.COUNTRY.BS,g:"1",index:27,h:!0},bt:{name:V.COUNTRY.BT,g:"975",index:146},bw:{name:V.COUNTRY.BW,g:"267",index:219},by:{name:V.COUNTRY.BY,g:"375",index:83},bz:{name:V.COUNTRY.BZ,g:"501",index:36},ca:{name:V.COUNTRY.CA,g:"1",index:106,
h:!0},cc:{name:V.COUNTRY.CC,g:"61",index:231,h:!0},cd:{name:V.COUNTRY.CD,g:"243",index:117},cf:{name:V.COUNTRY.CF,g:"236",index:145},cg:{name:V.COUNTRY.CG,g:"242",index:141},ch:{name:V.COUNTRY.CH,g:"41",index:101},ci:{name:V.COUNTRY.CI,g:"225",index:129},ck:{name:V.COUNTRY.CK,g:"682",index:183},cl:{name:V.COUNTRY.CL,g:"56",index:103},cm:{name:V.COUNTRY.CM,g:"237",index:165},cn:{name:V.COUNTRY.CN,g:"86",index:63},co:{name:V.COUNTRY.CO,g:"57",index:24},cr:{name:V.COUNTRY.CR,g:"506",index:168},cu:{name:V.COUNTRY.CU,
g:"53",index:58},cv:{name:V.COUNTRY.CV,g:"238",index:214},cw:{name:V.COUNTRY.CW,g:"599",index:221},cx:{name:V.COUNTRY.CX,g:"61",index:232,h:!0},cy:{name:V.COUNTRY.CY,g:"357",index:43},cz:{name:V.COUNTRY.CZ,g:"420",index:182},de:{name:V.COUNTRY.DE,g:"49",index:203},dj:{name:V.COUNTRY.DJ,g:"253",index:169},dk:{name:V.COUNTRY.DK,g:"45",index:107},dm:{name:V.COUNTRY.DM,g:"1",index:197,h:!0},"do":{name:V.COUNTRY.DO,g:"1",index:118,h:!0},dz:{name:V.COUNTRY.DZ,g:"213",index:40},ec:{name:V.COUNTRY.EC,g:"593",
index:90},ee:{name:V.COUNTRY.EE,g:"372",index:196},eg:{name:V.COUNTRY.EG,g:"20",index:178},eh:{name:V.COUNTRY.EH,g:"212",index:233,h:!0},er:{name:V.COUNTRY.ER,g:"291",index:55},es:{name:V.COUNTRY.ES,g:"34",index:87},et:{name:V.COUNTRY.ET,g:"251",index:198},fi:{name:V.COUNTRY.FI,g:"358",index:151},fj:{name:V.COUNTRY.FJ,g:"679",index:147},fk:{name:V.COUNTRY.FK,g:"500",index:224},fm:{name:V.COUNTRY.FM,g:"691",index:136},fo:{name:V.COUNTRY.FO,g:"298",index:84},fr:{name:V.COUNTRY.FR,g:"33",index:19},ga:{name:V.COUNTRY.GA,
g:"241",index:68},gb:{name:V.COUNTRY.GB,g:"44",index:5},gd:{name:V.COUNTRY.GD,g:"1",index:195,h:!0},ge:{name:V.COUNTRY.GE,g:"995",index:66},gf:{name:V.COUNTRY.GF,g:"594",index:19},gg:{name:V.COUNTRY.GG,g:"44",index:228,h:!0},gh:{name:V.COUNTRY.GH,g:"233",index:170},gi:{name:V.COUNTRY.GI,g:"350",index:20},gl:{name:V.COUNTRY.GL,g:"299",index:138},gm:{name:V.COUNTRY.GM,g:"220",index:48},gn:{name:V.COUNTRY.GN,g:"224",index:207},gp:{name:V.COUNTRY.GP,g:"590",index:30},gq:{name:V.COUNTRY.GQ,g:"240",index:116},
gr:{name:V.COUNTRY.GR,g:"30",index:11},gt:{name:V.COUNTRY.GT,g:"502",index:71},gu:{name:V.COUNTRY.GU,g:"1",index:192,h:!0},gw:{name:V.COUNTRY.GW,g:"245",index:153},gy:{name:V.COUNTRY.GY,g:"592",index:61},hk:{name:V.COUNTRY.HK,g:"852",index:218},hn:{name:V.COUNTRY.HN,g:"504",index:174},hr:{name:V.COUNTRY.HR,g:"385",index:69},ht:{name:V.COUNTRY.HT,g:"509",index:23},hu:{name:V.COUNTRY.HU,g:"36",index:53},id:{name:V.COUNTRY.ID,g:"62",index:156},ie:{name:V.COUNTRY.IE,g:"353",index:157},il:{name:V.COUNTRY.IL,
g:"972",index:25},im:{name:V.COUNTRY.IM,g:"44",index:229,h:!0},"in":{name:V.COUNTRY.IN,g:"91",index:132},io:{name:V.COUNTRY.IO,g:"246",index:5},iq:{name:V.COUNTRY.IQ,g:"964",index:50},ir:{name:V.COUNTRY.IR,g:"98",index:161},is:{name:V.COUNTRY.IS,g:"354",index:159},it:{name:V.COUNTRY.IT,g:"39",index:9},je:{name:V.COUNTRY.JE,g:"44",index:230,h:!0},jm:{name:V.COUNTRY.JM,g:"1",index:135,h:!0},jo:{name:V.COUNTRY.JO,g:"962",index:112},jp:{name:V.COUNTRY.JP,g:"81",index:31},ke:{name:V.COUNTRY.KE,g:"254",
index:212},kg:{name:V.COUNTRY.KG,g:"996",index:126},kh:{name:V.COUNTRY.KH,g:"855",index:17},ki:{name:V.COUNTRY.KI,g:"686",index:28},km:{name:V.COUNTRY.KM,g:"269",index:110},kn:{name:V.COUNTRY.KN,g:"1",index:6,h:!0},kp:{name:V.COUNTRY.KP,g:"850",index:142},kr:{name:V.COUNTRY.KR,g:"82",index:181},kw:{name:V.COUNTRY.KW,g:"965",index:202},ky:{name:V.COUNTRY.KY,g:"1",index:22,h:!0},kz:{name:V.COUNTRY.KZ,g:"7",index:92,h:!0},la:{name:V.COUNTRY.LA,g:"856",index:33},lb:{name:V.COUNTRY.LB,g:"961",index:95},
lc:{name:V.COUNTRY.LC,g:"1",index:108,h:!0},li:{name:V.COUNTRY.LI,g:"423",index:75},lk:{name:V.COUNTRY.LK,g:"94",index:213},lr:{name:V.COUNTRY.LR,g:"231",index:166},ls:{name:V.COUNTRY.LS,g:"266",index:177},lt:{name:V.COUNTRY.LT,g:"370",index:85},lu:{name:V.COUNTRY.LU,g:"352",index:113},lv:{name:V.COUNTRY.LV,g:"371",index:154},ly:{name:V.COUNTRY.LY,g:"218",index:8},ma:{name:V.COUNTRY.MA,g:"212",index:189},mc:{name:V.COUNTRY.MC,g:"377",index:70},md:{name:V.COUNTRY.MD,g:"373",index:217},me:{name:V.COUNTRY.ME,
g:"382",index:175},mf:{name:V.COUNTRY.MF,g:"590",index:5,h:!0},mg:{name:V.COUNTRY.MG,g:"261",index:98},mh:{name:V.COUNTRY.MH,g:"692",index:86},mk:{name:V.COUNTRY.MK,g:"389",index:104},ml:{name:V.COUNTRY.ML,g:"223",index:204},mm:{name:V.COUNTRY.MM,g:"95",index:1},mn:{name:V.COUNTRY.MN,g:"976",index:206},mo:{name:V.COUNTRY.MO,g:"853",index:209},mp:{name:V.COUNTRY.MP,g:"1",index:54,h:!0},mq:{name:V.COUNTRY.MQ,g:"596",index:14},mr:{name:V.COUNTRY.MR,g:"222",index:18},ms:{name:V.COUNTRY.MS,g:"1",index:44,
h:!0},mt:{name:V.COUNTRY.MT,g:"356",index:120},mu:{name:V.COUNTRY.MU,g:"230",index:176},mv:{name:V.COUNTRY.MV,g:"960",index:47},mw:{name:V.COUNTRY.MW,g:"265",index:173},mx:{name:V.COUNTRY.MX,g:"52",index:162},my:{name:V.COUNTRY.MY,g:"60",index:148},mz:{name:V.COUNTRY.MZ,g:"258",index:49},na:{name:V.COUNTRY.NA,g:"264",index:149},nc:{name:V.COUNTRY.NC,g:"687",index:97},ne:{name:V.COUNTRY.NE,g:"227",index:42},nf:{name:V.COUNTRY.NF,g:"672",index:15},ng:{name:V.COUNTRY.NG,g:"234",index:201},ni:{name:V.COUNTRY.NI,
g:"505",index:10},nl:{name:V.COUNTRY.NL,g:"31",index:111},no:{name:V.COUNTRY.NO,g:"47",index:64},np:{name:V.COUNTRY.NP,g:"977",index:7},nr:{name:V.COUNTRY.NR,g:"674",index:137},nu:{name:V.COUNTRY.NU,g:"683",index:167},nz:{name:V.COUNTRY.NZ,g:"64",index:119},om:{name:V.COUNTRY.OM,g:"968",index:199},pa:{name:V.COUNTRY.PA,g:"507",index:65},pe:{name:V.COUNTRY.PE,g:"51",index:72},pf:{name:V.COUNTRY.PF,g:"689",index:133},pg:{name:V.COUNTRY.PG,g:"675",index:114},ph:{name:V.COUNTRY.PH,g:"63",index:143},pk:{name:V.COUNTRY.PK,
g:"92",index:163},pl:{name:V.COUNTRY.PL,g:"48",index:89},pm:{name:V.COUNTRY.PM,g:"508",index:81},pr:{name:V.COUNTRY.PR,g:"1",index:35,h:!0},ps:{name:V.COUNTRY.PS,g:"970",index:91},pt:{name:V.COUNTRY.PT,g:"351",index:39},pw:{name:V.COUNTRY.PW,g:"680",index:16},py:{name:V.COUNTRY.PY,g:"595",index:190},qa:{name:V.COUNTRY.QA,g:"974",index:34},re:{name:V.COUNTRY.RE,g:"262",index:19},ro:{name:V.COUNTRY.RO,g:"40",index:52},rs:{name:V.COUNTRY.RS,g:"381",index:200},ru:{name:V.COUNTRY.RU,g:"7",index:51},rw:{name:V.COUNTRY.RW,
g:"250",index:216},sa:{name:V.COUNTRY.SA,g:"966",index:3},sb:{name:V.COUNTRY.SB,g:"677",index:80},sc:{name:V.COUNTRY.SC,g:"248",index:78},sd:{name:V.COUNTRY.SD,g:"249",index:26},se:{name:V.COUNTRY.SE,g:"46",index:29},sg:{name:V.COUNTRY.SG,g:"65",index:2},sh:{name:V.COUNTRY.SH,g:"290",index:37},si:{name:V.COUNTRY.SI,g:"386",index:93},sj:{name:V.COUNTRY.SJ,g:"47",index:64,h:!0},sk:{name:V.COUNTRY.SK,g:"421",index:179},sl:{name:V.COUNTRY.SL,g:"232",index:57},sm:{name:V.COUNTRY.SM,g:"378",index:171},
sn:{name:V.COUNTRY.SN,g:"221",index:172},so:{name:V.COUNTRY.SO,g:"252",index:105},sr:{name:V.COUNTRY.SR,g:"597",index:215},ss:{name:V.COUNTRY.SS,g:"211",index:222},st:{name:V.COUNTRY.ST,g:"239",index:194},sv:{name:V.COUNTRY.SV,g:"503",index:127},sx:{name:V.COUNTRY.SX,g:"1",index:225,h:!0},sy:{name:V.COUNTRY.SY,g:"963",index:144},sz:{name:V.COUNTRY.SZ,g:"268",index:184},ta:{name:V.COUNTRY.TA,g:"290",index:234,h:!0},tc:{name:V.COUNTRY.TC,g:"1",index:100,h:!0},td:{name:V.COUNTRY.TD,g:"235",index:62},
tg:{name:V.COUNTRY.TG,g:"228",index:46},th:{name:V.COUNTRY.TH,g:"66",index:73},tj:{name:V.COUNTRY.TJ,g:"992",index:13},tk:{name:V.COUNTRY.TK,g:"690",index:223},tl:{name:V.COUNTRY.TL,g:"670",index:226},tm:{name:V.COUNTRY.TM,g:"993",index:205},tn:{name:V.COUNTRY.TN,g:"216",index:41},to:{name:V.COUNTRY.TO,g:"676",index:82},tr:{name:V.COUNTRY.TR,g:"90",index:125},tt:{name:V.COUNTRY.TT,g:"1",index:32,h:!0},tv:{name:V.COUNTRY.TV,g:"688",index:21},tw:{name:V.COUNTRY.TW,g:"886",index:38},tz:{name:V.COUNTRY.TZ,
g:"255",index:185},ua:{name:V.COUNTRY.UA,g:"380",index:160},ug:{name:V.COUNTRY.UG,g:"256",index:88},us:{name:V.COUNTRY.US,g:"1",index:4},uy:{name:V.COUNTRY.UY,g:"598",index:210},uz:{name:V.COUNTRY.UZ,g:"998",index:76},va:{name:V.COUNTRY.VA,g:"39",index:188,h:!0},vc:{name:V.COUNTRY.VC,g:"1",index:211,h:!0},ve:{name:V.COUNTRY.VE,g:"58",index:79},vg:{name:V.COUNTRY.VG,g:"1",index:109,h:!0},vi:{name:V.COUNTRY.VI,g:"1",index:140,h:!0},vn:{name:V.COUNTRY.VN,g:"84",index:74},vu:{name:V.COUNTRY.VU,g:"678",
index:96},wf:{name:V.COUNTRY.WF,g:"681",index:19},ws:{name:V.COUNTRY.WS,g:"685",index:186},xk:{name:V.COUNTRY.XK,g:"383",index:227},ye:{name:V.COUNTRY.YE,g:"967",index:130},yt:{name:V.COUNTRY.YT,g:"262",index:19,h:!0},za:{name:V.COUNTRY.ZA,g:"27",index:191},zm:{name:V.COUNTRY.ZM,g:"260",index:124},zw:{name:V.COUNTRY.ZW,g:"263",index:164}};var W=function(){y.apply(this,arguments)};v(W,y);
W.prototype.l=function(){var b=this.i.querySelector("SELECT".toString()),c=document.createDocumentFragment(),d=Object.keys(pa),e=(this.i.dataset.regionCode||"").toLowerCase();d=w(d);for(var f=d.next();!f.done;f=d.next()){var g=f.value;f=pa[g];var k=f.g,n=f.name;f=g.toLowerCase()===e;var t=document.createElement("OPTION".toString());t.value=g;g="(+"+k+") "+n;g instanceof M||(g=String(g).replace(/&/g,"&amp;").replace(/</g,"&lt;").replace(/>/g,"&gt;").replace(/"/g,"&quot;").replace(/'/g,"&apos;"),I===
void 0&&(I=ha()),k=I,g=new M(k?k.createHTML(g):g));t.textContent=g.toString();f&&(t.selected=!0);c.appendChild(t)}b.appendChild(c)};var X=function(){y.apply(this,arguments)};v(X,y);X.prototype.l=function(){var b=this;this.m=[].concat(ea(this.i.querySelectorAll('input[type="checkbox"]:not(input[type="checkbox"][data-is-select-all])')));if(this.j=this.i.querySelector('input[type="checkbox"][data-is-select-all]'))qa(this),this.i.addEventListener("change",function(c){c.target&&(c=c.target,c.type==="checkbox"&&(c===b.j?ra(b,c.checked):qa(b)))})};
var ra=function(b,c){b.m.forEach(function(d){d.checked=c})},qa=function(b){var c=b.m.filter(function(d){return d.checked}).length;c===0?(b.j.indeterminate=!1,b.j.checked=!1):c>0&&c<b.m.length?(b.j.indeterminate=!0,b.j.checked=!0):c===b.m.length&&(b.j.indeterminate=!1,b.j.checked=!0)};P("AccountChooser",C);P("CaptchaInput",Q);P("Card",E);P("CountrySelect",W);P("EmailInput",R);P("Footer",N);P("IdentifierInput",U);P("RecaptchaInput",T);P("SelectionInput",X);for(var sa=[],ta=w([].slice.call(document.querySelectorAll("[data-auto-init]"))),Y=ta.next();!Y.done;Y=ta.next()){var Z=Y.value,ua=Z.getAttribute("data-auto-init");if(!ua)throw Error("auto-init attribute requires a value.");var va=new O[ua](Z);sa.push(va);Z.removeAttribute("data-auto-init")};}).call(this);
</script></div></div></body>